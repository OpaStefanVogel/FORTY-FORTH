library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity FortyForthProcessor is
  Port (
    CLK_I: in STD_LOGIC;
    DAT_I: in STD_LOGIC_VECTOR (15 downto 0);
    ADR_O: out STD_LOGIC_VECTOR (15 downto 0);
    DAT_O: out STD_LOGIC_VECTOR (15 downto 0);
    WE_O: out STD_LOGIC;
    
    -- EMIT --
    EMIT_ABGESCHICKT: out STD_LOGIC;
    EMIT_BYTE: out STD_LOGIC_VECTOR (7 downto 0);
    EMIT_ANGEKOMMEN: in STD_LOGIC;
    
     -- EMIT --
    KEY_ABGESCHICKT: in STD_LOGIC;
    KEY_BYTE: in STD_LOGIC_VECTOR (7 downto 0);
    KEY_ANGEKOMMEN: out STD_LOGIC;

   -- nur zur Simulation und Fehlersuche:
    PC_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    PD_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    SP_SIM: out integer;
    A_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    B_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    C_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    D_SIM: out STD_LOGIC_VECTOR (15 downto 0)
    );
end FortyForthProcessor;

architecture Step_9 of FortyForthProcessor is

constant SHA: STD_LOGIC_VECTOR (10*16-1 downto 0):=
  x"b2cc26074b713be1a669ef7cb895d72533c8dad9";
type REG is array(0 to 3) of STD_LOGIC_VECTOR (15 downto 0);
type RAMTYPE is array(0 to 8*1024-1) of STD_LOGIC_VECTOR (15 downto 0);
-- Programmspeicher 0000H-1FFFH
signal ProgRAM: RAMTYPE:=(
-- 
  x"4010",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 0000-000F 
  x"476D",x"A003",x"44BA",x"9001",x"A003",x"B300",x"8000",x"8FFA",x"0000",x"11A4",x"0000",x"0000",x"0000",x"0000",x"1199",x"118F", -- 0010-001F 
  x"4000",x"A003",x"4000",x"A003",x"4000",x"A003",x"448B",x"A003",x"0000",x"3000",x"0001",x"4780",x"0029",x"45F2",x"B200",x"A003", -- 0020-002F 
  x"FFF8",x"3002",x"0001",x"4780",x"0000",x"2F10",x"A009",x"A003",x"FFF8",x"3004",x"0001",x"478E",x"0001",x"2F10",x"A009",x"A003", -- 0030-003F 
  x"FFF8",x"3006",x"0007",x"4780",x"0020",x"45F2",x"466C",x"46AC",x"B300",x"46B5",x"A003",x"FFF5",x"300E",x"0006",x"4787",x"42D4", -- 0040-004F 
  x"B501",x"4287",x"42E7",x"A00A",x"A003",x"FFF6",x"3015",x"0004",x"478E",x"51EF",x"A003",x"42AE",x"B502",x"C000",x"429C",x"A00E", -- 0050-005F 
  x"9001",x"404E",x"4307",x"A003",x"FFF1",x"301A",x"000B",x"4787",x"42D4",x"A00A",x"2F10",x"A00A",x"9001",x"4059",x"A003",x"FFF5", -- 0060-006F 
  x"3026",x"0008",x"478E",x"46BE",x"4067",x"4307",x"4778",x"A003",x"FFF7",x"302F",x"0006",x"4068",x"2800",x"FFFB",x"3036",x"0002", -- 0070-007F 
  x"4068",x"2801",x"FFFB",x"3039",x"0002",x"4068",x"2802",x"FFFB",x"303C",x"0002",x"4068",x"2803",x"FFFB",x"303F",x"0004",x"4068", -- 0080-008F 
  x"2F00",x"FFFB",x"3044",x"0009",x"4068",x"2F01",x"FFFB",x"304E",x"0003",x"4068",x"2F02",x"FFFB",x"3052",x"0007",x"4068",x"2F03", -- 0090-009F 
  x"FFFB",x"305A",x"0007",x"4068",x"2F04",x"FFFB",x"3062",x"0004",x"4068",x"2F05",x"FFFB",x"3067",x"0007",x"4068",x"2F06",x"FFFB", -- 00A0-00AF 
  x"306F",x"0004",x"4068",x"2F07",x"FFFB",x"3074",x"0004",x"4068",x"2F08",x"FFFB",x"3079",x"0003",x"4068",x"2F09",x"FFFB",x"307D", -- 00B0-00BF 
  x"0003",x"4068",x"2F0A",x"FFFB",x"3081",x"0003",x"4068",x"2F0B",x"FFFB",x"3085",x"0003",x"4068",x"2F0C",x"FFFB",x"3089",x"0003", -- 00C0-00CF 
  x"4068",x"2F0D",x"FFFB",x"308D",x"0007",x"4068",x"2F0E",x"FFFB",x"3095",x"0002",x"4068",x"2F0F",x"FFFB",x"3098",x"0004",x"4068", -- 00D0-00DF 
  x"2F10",x"FFFB",x"309D",x"0003",x"4068",x"2F11",x"FFFB",x"30A1",x"0004",x"4068",x"2F12",x"FFFB",x"30A6",x"0005",x"4068",x"2F13", -- 00E0-00EF 
  x"FFFB",x"30AC",x"0006",x"4068",x"2F14",x"FFFB",x"30B3",x"0003",x"4068",x"2F15",x"FFFB",x"30B7",x"0009",x"4068",x"2F16",x"FFFB", -- 00F0-00FF 
  x"30C1",x"000C",x"4068",x"2F17",x"FFFB",x"30CE",x"0007",x"4068",x"01B2",x"FFFB",x"30D6",x"0006",x"4068",x"A003",x"FFFB",x"30DD", -- 0100-010F 
  x"0008",x"4787",x"42D4",x"2F10",x"A00A",x"9003",x"A00A",x"4307",x"8001",x"4312",x"A003",x"FFF3",x"30E6",x"0005",x"478E",x"46BE", -- 0110-011F 
  x"4111",x"4307",x"404F",x"A003",x"4307",x"4778",x"A003",x"FFF4",x"30EC",x"0005",x"4112",x"A000",x"A003",x"FFFA",x"30F2",x"0002", -- 0120-012F 
  x"4112",x"A001",x"A003",x"FFFA",x"30F5",x"0002",x"4112",x"A002",x"A003",x"FFFA",x"30F8",x"0002",x"4112",x"A00D",x"A003",x"FFFA", -- 0130-013F 
  x"30FB",x"0003",x"4112",x"A00F",x"A003",x"FFFA",x"30FF",x"0008",x"4112",x"A005",x"A003",x"FFFA",x"3108",x"0003",x"4112",x"A00B", -- 0140-014F 
  x"A003",x"FFFA",x"310C",x"0003",x"4112",x"A008",x"A003",x"FFFA",x"3110",x"0002",x"4112",x"A00E",x"A003",x"FFFA",x"3113",x"0007", -- 0150-015F 
  x"4112",x"A00C",x"A003",x"FFFA",x"311B",x"0001",x"4112",x"A007",x"A003",x"FFFA",x"311D",x"0001",x"4112",x"A009",x"A003",x"FFFA", -- 0160-016F 
  x"311F",x"0001",x"4112",x"A00A",x"A003",x"FFFA",x"3121",x"0004",x"4112",x"B412",x"A003",x"FFFA",x"3126",x"0004",x"4112",x"B502", -- 0170-017F 
  x"A003",x"FFFA",x"312B",x"0003",x"4112",x"B501",x"A003",x"FFFA",x"312F",x"0003",x"4112",x"B434",x"A003",x"FFFA",x"3133",x"0004", -- 0180-018F 
  x"4112",x"B300",x"A003",x"FFFA",x"3138",x"0005",x"4112",x"B43C",x"A003",x"FFFA",x"313E",x"0005",x"4112",x"B60C",x"A003",x"FFFA", -- 0190-019F 
  x"3144",x"0004",x"4112",x"B603",x"A003",x"FFFA",x"3149",x"0005",x"4112",x"B200",x"A003",x"FFFA",x"314F",x"0004",x"4112",x"8000", -- 01A0-01AF 
  x"A003",x"FFFA",x"3154",x"0002",x"478E",x"2F13",x"A00A",x"A009",x"0001",x"2F13",x"42C9",x"A003",x"FFF5",x"3157",x"0002",x"478E", -- 01B0-01BF 
  x"2F13",x"A00A",x"4059",x"B501",x"4307",x"B412",x"B501",x"A00A",x"41B5",x"4287",x"B412",x"0001",x"428E",x"B501",x"A00D",x"9FF5", -- 01C0-01CF 
  x"B200",x"0020",x"41B5",x"A003",x"FFE8",x"315A",x"0007",x"4787",x"45F2",x"2F10",x"A00A",x"9003",x"41C0",x"42D4",x"46B5",x"A003", -- 01D0-01DF 
  x"FFF4",x"3162",x"0005",x"478E",x"46BE",x"0001",x"2F10",x"A009",x"4307",x"41D7",x"FFFF",x"2F15",x"42C9",x"A003",x"FFF2",x"3168", -- 01E0-01EF 
  x"0001",x"0022",x"41D8",x"A003",x"FFFA",x"316A",x"0002",x"0022",x"41D8",x"433F",x"A003",x"FFF9",x"316D",x"0004",x"478E",x"2F0F", -- 01F0-01FF 
  x"A00A",x"A003",x"FFF9",x"3172",x"0005",x"478E",x"0008",x"A003",x"FFFA",x"3178",x"0006",x"478E",x"0009",x"A003",x"FFFA",x"317F", -- 0200-020F 
  x"0006",x"478E",x"1000",x"42B5",x"B412",x"0FFF",x"A008",x"A00E",x"A003",x"FFF5",x"3186",x"0005",x"478E",x"2F0F",x"42C9",x"A003", -- 0210-021F 
  x"FFF9",x"318C",x"0007",x"478E",x"41FF",x"4287",x"428E",x"4206",x"4212",x"4307",x"A003",x"FFF5",x"3194",x"0008",x"478E",x"41FF", -- 0220-022F 
  x"4287",x"428E",x"420C",x"4212",x"4307",x"A003",x"FFF5",x"319D",x"0005",x"4780",x"41FF",x"A003",x"FFFA",x"31A3",x"0005",x"4780", -- 0230-023F 
  x"4224",x"A003",x"FFFA",x"31A9",x"0005",x"4780",x"422F",x"A003",x"FFFA",x"31AF",x"0002",x"4780",x"420C",x"0001",x"421D",x"41FF", -- 0240-024F 
  x"A003",x"FFF7",x"31B2",x"0006",x"4780",x"41FF",x"B502",x"428E",x"B434",x"4212",x"B412",x"0001",x"428E",x"A009",x"A003",x"FFF2", -- 0250-025F 
  x"31B9",x"0004",x"4780",x"0001",x"421D",x"4254",x"4206",x"41FF",x"A003",x"FFF6",x"31BE",x"0005",x"4780",x"424B",x"A003",x"FFFA", -- 0260-026F 
  x"31C4",x"0006",x"4780",x"B434",x"423F",x"4254",x"A003",x"FFF8",x"31CB",x"0002",x"478E",x"A00A",x"A003",x"FFFA",x"31CE",x"0002", -- 0270-027F 
  x"478E",x"A009",x"A003",x"FFFA",x"31D1",x"0002",x"478E",x"0001",x"A007",x"A003",x"FFF9",x"31D4",x"0001",x"478E",x"A000",x"A007", -- 0280-028F 
  x"A003",x"FFF9",x"31D6",x"0001",x"478E",x"428E",x"A00D",x"A003",x"FFF9",x"31D8",x"0002",x"478E",x"404F",x"8000",x"A007",x"B412", -- 0290-029F 
  x"A00B",x"404F",x"8000",x"A007",x"0000",x"A001",x"B300",x"A00D",x"A00B",x"A003",x"FFEE",x"31DB",x"0001",x"478E",x"B412",x"429C", -- 02A0-02AF 
  x"A003",x"FFF9",x"31DD",x"0001",x"478E",x"0000",x"B434",x"B434",x"A002",x"B412",x"B300",x"A003",x"FFF5",x"31DF",x"0003",x"478E", -- 02B0-02BF 
  x"31E3",x"0004",x"41F9",x"8FFC",x"A003",x"FFF7",x"31E8",x"0002",x"478E",x"B412",x"B502",x"A00A",x"A007",x"B412",x"A009",x"A003", -- 02C0-02CF 
  x"FFF5",x"31EB",x"0002",x"478E",x"2802",x"A00A",x"4287",x"A00A",x"2802",x"A00A",x"4287",x"2802",x"B603",x"A00A",x"A00A",x"B412", -- 02D0-02DF 
  x"A009",x"A009",x"A003",x"FFED",x"31EE",x"0002",x"478E",x"2802",x"A00A",x"B501",x"FFFF",x"A007",x"2802",x"B603",x"A00A",x"A00A", -- 02E0-02EF 
  x"B412",x"B501",x"FFFF",x"A007",x"2802",x"A009",x"A009",x"A009",x"A009",x"A003",x"FFE9",x"31F1",x"0001",x"478E",x"2802",x"A00A", -- 02F0-02FF 
  x"4287",x"A00A",x"A003",x"FFF7",x"31F3",x"0001",x"478E",x"2F0F",x"A00A",x"A009",x"0001",x"2F0F",x"42C9",x"A003",x"FFF5",x"31F5", -- 0300-030F 
  x"0007",x"478E",x"2803",x"A009",x"A003",x"FFF9",x"31FD",x"0003",x"478E",x"0012",x"4312",x"A003",x"FFF9",x"3201",x"0004",x"478E", -- 0310-031F 
  x"0149",x"4312",x"A003",x"FFF9",x"3206",x"0005",x"478E",x"0000",x"B412",x"0010",x"A002",x"B412",x"A003",x"FFF6",x"320C",x"0003", -- 0320-032F 
  x"478E",x"B501",x"000A",x"429C",x"9001",x"8002",x"0007",x"A007",x"0030",x"A007",x"A003",x"FFF2",x"3210",x"0004",x"478E",x"B501", -- 0330-033F 
  x"9009",x"B412",x"B501",x"427B",x"4320",x"4287",x"B412",x"0001",x"428E",x"8FF5",x"B200",x"A003",x"FFEF",x"3215",x"0003",x"478E", -- 0340-034F 
  x"4327",x"4331",x"4320",x"4327",x"4331",x"4320",x"4327",x"4331",x"4320",x"4327",x"4331",x"4320",x"B300",x"A003",x"FFEE",x"3219", -- 0350-035F 
  x"0002",x"478E",x"4350",x"0020",x"4320",x"A003",x"FFF8",x"321C",x"0001",x"478E",x"4362",x"A003",x"FFFA",x"321E",x"0001",x"478E", -- 0360-036F 
  x"A00A",x"436A",x"A003",x"FFF9",x"3220",x"0002",x"478E",x"2F07",x"A00A",x"2F0F",x"A00A",x"428E",x"2F10",x"A00A",x"A00D",x"A00B", -- 0370-037F 
  x"A00E",x"2F00",x"A00A",x"A00D",x"A00B",x"A008",x"9028",x"003C",x"4320",x"3223",x"0003",x"41F9",x"2F07",x"A00A",x"436A",x"2F06", -- 0380-038F 
  x"A00A",x"436A",x"003C",x"4320",x"3227",x"0004",x"41F9",x"003C",x"4320",x"322C",x"0003",x"41F9",x"2F0F",x"A00A",x"436A",x"2F13", -- 0390-039F 
  x"A00A",x"436A",x"003C",x"4320",x"3230",x"0004",x"41F9",x"2F0F",x"A00A",x"2F07",x"A009",x"2F13",x"A00A",x"2F06",x"A009",x"000A", -- 03A0-03AF 
  x"4320",x"A003",x"FFC1",x"3235",x"000A",x"478E",x"A003",x"FFFB",x"3240",x"0007",x"478E",x"4377",x"3248",x"0019",x"41F9",x"0020", -- 03B0-03BF 
  x"4320",x"0008",x"4320",x"4319",x"001B",x"4295",x"9FF8",x"A003",x"FFEF",x"3262",x"0005",x"478E",x"B501",x"2F0E",x"A009",x"0000", -- 03C0-03CF 
  x"2F10",x"A009",x"4377",x"2F0A",x"A00A",x"2F0C",x"A00A",x"2F0A",x"A00A",x"428E",x"0001",x"428E",x"433F",x"3268",x"0003",x"41F9", -- 03D0-03DF 
  x"326C",x"000A",x"41F3",x"46D3",x"4377",x"3277",x"0016",x"41F9",x"436A",x"43BB",x"4720",x"A003",x"FFDC",x"328E",x"0004",x"478E", -- 03E0-03EF 
  x"2801",x"A00A",x"2F15",x"A009",x"A003",x"FFF7",x"3293",x"0004",x"478E",x"2801",x"A00A",x"2F15",x"A00A",x"428E",x"9002",x"0009", -- 03F0-03FF 
  x"43CC",x"A003",x"FFF3",x"3298",x"0005",x"478E",x"0001",x"A007",x"2F17",x"A00A",x"B502",x"428E",x"B501",x"2F17",x"A009",x"A009", -- 0400-040F 
  x"A003",x"FFF1",x"329E",x"0009",x"478E",x"2F17",x"A00A",x"B501",x"A00A",x"A007",x"2F17",x"A009",x"A003",x"FFF4",x"32A8",x"0002", -- 0410-041F 
  x"478E",x"2F17",x"A00A",x"0001",x"A007",x"A003",x"FFF7",x"32AB",x"0002",x"478E",x"2F17",x"A00A",x"0002",x"A007",x"A003",x"FFF7", -- 0420-042F 
  x"32AE",x"0002",x"478E",x"2F17",x"A00A",x"0003",x"A007",x"A003",x"FFF7",x"32B1",x"0002",x"478E",x"2F17",x"A00A",x"0004",x"A007", -- 0430-043F 
  x"A003",x"FFF7",x"32B4",x"0002",x"478E",x"2F17",x"A00A",x"0005",x"A007",x"A003",x"FFF7",x"32B7",x"0002",x"478E",x"2F17",x"A00A", -- 0440-044F 
  x"0006",x"A007",x"A003",x"FFF7",x"32BA",x"0002",x"478E",x"2F17",x"A00A",x"0007",x"A007",x"A003",x"FFF7",x"32BD",x"0002",x"478E", -- 0450-045F 
  x"2F17",x"A00A",x"0008",x"A007",x"A003",x"FFF7",x"32C0",x"0001",x"4780",x"0020",x"45F2",x"466C",x"46AC",x"B300",x"4287",x"2F10", -- 0460-046F 
  x"A00A",x"9001",x"4059",x"A003",x"FFF1",x"32C2",x"0005",x"478E",x"B501",x"A00A",x"0001",x"A007",x"B501",x"03FF",x"A008",x"0000", -- 0470-047F 
  x"4295",x"9002",x"0400",x"428E",x"B412",x"A009",x"A003",x"FFED",x"32C8",x"0007",x"478E",x"2800",x"A00A",x"B501",x"0008",x"429C", -- 0480-048F 
  x"9009",x"0018",x"A007",x"A00A",x"B501",x"9002",x"B501",x"4312",x"B300",x"8018",x"2F03",x"A00A",x"A009",x"2F03",x"4478",x"2F03", -- 0490-049F 
  x"A00A",x"2F04",x"A00A",x"428E",x"03FF",x"A008",x"0080",x"42AE",x"9009",x"2F05",x"A00A",x"A00D",x"9005",x"FFFF",x"2F05",x"A009", -- 04A0-04AF 
  x"0013",x"4320",x"0000",x"2800",x"A009",x"A003",x"FFD1",x"32D0",x"0008",x"478E",x"2F04",x"A00A",x"2F03",x"A00A",x"4295",x"9003", -- 04B0-04BF 
  x"0000",x"0000",x"8018",x"2F04",x"A00A",x"A00A",x"FFFF",x"2F04",x"4478",x"2F03",x"A00A",x"2F04",x"A00A",x"428E",x"03FF",x"A008", -- 04C0-04CF 
  x"0020",x"429C",x"9008",x"2F05",x"A00A",x"9005",x"0000",x"2F05",x"A009",x"0011",x"4320",x"A003",x"FFDA",x"32D9",x"0006",x"478E", -- 04D0-04DF 
  x"0005",x"4406",x"4433",x"A009",x"442A",x"A009",x"442A",x"A00A",x"4445",x"A009",x"4319",x"B501",x"0014",x"4295",x"9004",x"B300", -- 04E0-04EF 
  x"442A",x"A00A",x"427B",x"B501",x"007F",x"4295",x"9002",x"B300",x"0008",x"B501",x"0008",x"4295",x"9012",x"4445",x"A00A",x"442A", -- 04F0-04FF 
  x"A00A",x"429C",x"900C",x"FFFF",x"442A",x"42C9",x"0001",x"4433",x"42C9",x"0008",x"4320",x"0020",x"4320",x"0008",x"4320",x"B501", -- 0500-050F 
  x"0020",x"429C",x"9001",x"8012",x"FFFF",x"4433",x"42C9",x"4433",x"A00A",x"A00F",x"9002",x"0006",x"43CC",x"B501",x"4320",x"B501", -- 0510-051F 
  x"442A",x"A00A",x"4281",x"0001",x"442A",x"42C9",x"B501",x"0020",x"429C",x"B502",x"0008",x"4295",x"A00B",x"A008",x"B412",x"001B", -- 0520-052F 
  x"4295",x"A00B",x"A008",x"4433",x"A00A",x"A00D",x"A00E",x"9FB2",x"0020",x"4320",x"4445",x"A00A",x"442A",x"A00A",x"4445",x"A00A", -- 0530-053F 
  x"428E",x"B603",x"A007",x"0000",x"B412",x"4281",x"4415",x"A003",x"FF94",x"32E0",x"0005",x"478E",x"B501",x"0030",x"429C",x"A00B", -- 0540-054F 
  x"B502",x"003A",x"429C",x"A008",x"B502",x"0041",x"429C",x"A00B",x"A00E",x"B501",x"9015",x"B412",x"0030",x"428E",x"B501",x"000A", -- 0550-055F 
  x"429C",x"A00B",x"9002",x"0007",x"428E",x"B501",x"2F08",x"A00A",x"429C",x"A00B",x"9004",x"B300",x"B300",x"0000",x"0000",x"B412", -- 0560-056F 
  x"A003",x"FFD7",x"32E6",x"0006",x"478E",x"51F1",x"A003",x"442A",x"A009",x"4421",x"A009",x"0000",x"442A",x"A00A",x"9063",x"B501", -- 0570-057F 
  x"4433",x"A009",x"0001",x"444E",x"A009",x"FFFF",x"4457",x"A009",x"4421",x"A00A",x"4433",x"A00A",x"A007",x"427B",x"002B",x"4295", -- 0580-058F 
  x"9009",x"4433",x"A00A",x"4287",x"4433",x"A009",x"0000",x"4457",x"A009",x"8016",x"4421",x"A00A",x"4433",x"A00A",x"A007",x"427B", -- 0590-059F 
  x"002D",x"4295",x"900D",x"4433",x"A00A",x"4287",x"4433",x"A009",x"0000",x"4457",x"A009",x"444E",x"A00A",x"A000",x"444E",x"A009", -- 05A0-05AF 
  x"4457",x"A00A",x"9FD2",x"4433",x"A00A",x"442A",x"A00A",x"429C",x"9029",x"4421",x"A00A",x"4433",x"A00A",x"A007",x"427B",x"B501", -- 05B0-05BF 
  x"9015",x"454C",x"A00B",x"9007",x"B300",x"442A",x"A00A",x"A000",x"442A",x"A009",x"800A",x"B412",x"2F08",x"A00A",x"42B5",x"A007", -- 05C0-05CF 
  x"4433",x"A00A",x"4287",x"4433",x"A009",x"8005",x"B300",x"4433",x"A00A",x"442A",x"A009",x"4433",x"A00A",x"442A",x"A00A",x"429C", -- 05D0-05DF 
  x"A00B",x"9FD7",x"444E",x"A00A",x"A00F",x"9001",x"A000",x"4433",x"A00A",x"442A",x"A00A",x"428E",x"4415",x"A003",x"FF83",x"32ED", -- 05E0-05EF 
  x"0004",x"478E",x"42E7",x"2F0C",x"A00A",x"2F0B",x"A009",x"2F0C",x"A00A",x"427B",x"42FE",x"4295",x"2F0C",x"A00A",x"2F0D",x"A00A", -- 05F0-05FF 
  x"429C",x"A008",x"9004",x"0001",x"2F0C",x"42C9",x"8FF0",x"2F0C",x"A00A",x"2F0B",x"A009",x"2F0C",x"A00A",x"427B",x"003C",x"4295", -- 0600-060F 
  x"9004",x"2F0C",x"A00A",x"2F0D",x"A009",x"2F0C",x"A00A",x"427B",x"42FE",x"4295",x"A00B",x"2F0C",x"A00A",x"2F0D",x"A00A",x"429C", -- 0610-061F 
  x"A008",x"9004",x"0001",x"2F0C",x"42C9",x"8FE5",x"2F0B",x"A00A",x"2F0C",x"A00A",x"B502",x"428E",x"B501",x"9003",x"0001",x"2F0C", -- 0620-062F 
  x"42C9",x"42D4",x"B300",x"A003",x"FFBA",x"32F2",x"0002",x"478E",x"42E7",x"B502",x"42FE",x"428E",x"9007",x"42D4",x"B300",x"B300", -- 0630-063F 
  x"B300",x"B300",x"0000",x"8023",x"42D4",x"B300",x"B412",x"0000",x"B603",x"428E",x"9016",x"42E7",x"42E7",x"B502",x"427B",x"B502", -- 0640-064F 
  x"427B",x"428E",x"9004",x"B300",x"B300",x"0000",x"0000",x"B501",x"9004",x"4287",x"B412",x"4287",x"B412",x"42D4",x"42D4",x"4287", -- 0650-065F 
  x"8FE7",x"B200",x"B300",x"9002",x"FFFF",x"8001",x"0000",x"A003",x"FFCC",x"32F5",x"0004",x"478E",x"42E7",x"42E7",x"0000",x"2F11", -- 0660-066F 
  x"A00A",x"2F01",x"A00A",x"9003",x"B501",x"A00A",x"A007",x"B501",x"4287",x"B501",x"A00A",x"B412",x"4287",x"A00A",x"42D4",x"42D4", -- 0670-067F 
  x"B603",x"42E7",x"42E7",x"4638",x"9003",x"B412",x"A00D",x"B412",x"B502",x"A00D",x"B502",x"A00A",x"A00D",x"A00B",x"A008",x"B502", -- 0680-068F 
  x"B501",x"A00A",x"A007",x"2F11",x"A00A",x"4295",x"A00B",x"A008",x"9004",x"B501",x"A00A",x"A007",x"8FDA",x"42D4",x"B300",x"42D4", -- 0690-069F 
  x"B434",x"A00D",x"9004",x"B300",x"B300",x"0000",x"0000",x"A003",x"FFC0",x"32FA",x"0004",x"478E",x"B412",x"0003",x"A007",x"B412", -- 06A0-06AF 
  x"A003",x"FFF7",x"32FF",x"0008",x"478E",x"404F",x"4000",x"A007",x"4307",x"A003",x"FFF7",x"3308",x"0006",x"478E",x"43F0",x"2F0F", -- 06B0-06BF 
  x"A00A",x"2F11",x"A00A",x"B502",x"428E",x"4307",x"2F11",x"A009",x"0020",x"45F2",x"41C0",x"0001",x"2F01",x"A009",x"A003",x"FFEB", -- 06C0-06CF 
  x"330F",x"0009",x"478E",x"2F0A",x"A00A",x"42E7",x"2F0B",x"A00A",x"42E7",x"2F0C",x"A00A",x"42E7",x"2F0D",x"A00A",x"42E7",x"B502", -- 06D0-06DF 
  x"A007",x"2F0D",x"A009",x"B501",x"2F0A",x"A009",x"B501",x"2F0B",x"A009",x"2F0C",x"A009",x"0020",x"45F2",x"B501",x"901F",x"B603", -- 06E0-06EF 
  x"466C",x"B501",x"9009",x"42E7",x"42E7",x"B200",x"42D4",x"42D4",x"46AC",x"B300",x"4312",x"8011",x"B200",x"B603",x"4575",x"9005", -- 06F0-06FF 
  x"B200",x"B300",x"0003",x"43CC",x"8008",x"B434",x"B300",x"B412",x"B300",x"2F10",x"A00A",x"9001",x"4059",x"8FDD",x"B200",x"42D4", -- 0700-070F 
  x"2F0D",x"A009",x"42D4",x"2F0C",x"A009",x"42D4",x"2F0B",x"A009",x"42D4",x"2F0A",x"A009",x"A003",x"FFB3",x"3319",x"0004",x"478E", -- 0710-071F 
  x"2F02",x"A00A",x"2802",x"A009",x"2F00",x"A00A",x"9006",x"003C",x"4320",x"331E",x"0004",x"41F9",x"8003",x"3323",x"0002",x"41F9", -- 0720-072F 
  x"4377",x"2F09",x"A00A",x"0100",x"44E0",x"B502",x"A00A",x"003C",x"4295",x"9002",x"B200",x"802B",x"2F00",x"A00A",x"900C",x"003C", -- 0730-073F 
  x"4320",x"3326",x"0003",x"41F9",x"46D3",x"003C",x"4320",x"332A",x"0004",x"41F9",x"801C",x"001B",x"4320",x"005B",x"4320",x"0033", -- 0740-074F 
  x"4320",x"0036",x"4320",x"006D",x"4320",x"46D3",x"2F10",x"A00A",x"A00D",x"9003",x"332F",x"0002",x"41F9",x"001B",x"4320",x"005B", -- 0750-075F 
  x"4320",x"0033",x"4320",x"0039",x"4320",x"006D",x"4320",x"8FC8",x"A003",x"FFB3",x"3332",x"0005",x"478E",x"3338",x"000B",x"41F9", -- 0760-076F 
  x"4377",x"4377",x"4720",x"A003",x"FFF5",x"3344",x"0006",x"478E",x"0000",x"2F01",x"A009",x"A003",x"FFF8",x"334B",x"000C",x"478E", -- 0770-077F 
  x"42D4",x"42E7",x"A003",x"FFF9",x"3358",x"000A",x"478E",x"42D4",x"46B5",x"A003",x"FFF9",x"3363",x"0003",x"478E",x"42D4",x"2F10", -- 0780-078F 
  x"A00A",x"9002",x"46B5",x"8001",x"42E7",x"A003",x"FFF4",x"3367",x"000A",x"478E",x"46BE",x"0001",x"2F10",x"A009",x"477F",x"A003", -- 0790-079F 
  x"FFF6",x"3372",x"0008",x"478E",x"46BE",x"0001",x"2F10",x"A009",x"4786",x"A003",x"FFF6",x"337B",x"0001",x"478E",x"46BE",x"0001", -- 07A0-07AF 
  x"2F10",x"A009",x"478D",x"A003",x"FFF6",x"337D",x"0001",x"4780",x"0000",x"2F10",x"A009",x"43F9",x"404F",x"A003",x"4307",x"4778", -- 07B0-07BF 
  x"A003",x"FFF3",x"337F",x"0005",x"478E",x"41FF",x"A003",x"FFFA",x"3385",x"0003",x"478E",x"47C5",x"A00A",x"9005",x"4327",x"B300", -- 07C0-07CF 
  x"4327",x"B300",x"8006",x"4327",x"4331",x"4320",x"4327",x"4331",x"4320",x"4327",x"4331",x"4320",x"4327",x"4331",x"4320",x"B300", -- 07D0-07DF 
  x"A003",x"FFE6",x"3389",x"0003",x"478E",x"338D",x"0001",x"41F9",x"0022",x"4320",x"47CB",x"0022",x"4320",x"338F",x"0001",x"41F9", -- 07E0-07EF 
  x"A003",x"FFF0",x"3391",x"0005",x"478E",x"47C5",x"A009",x"2F00",x"A00A",x"42E7",x"0000",x"2F00",x"A009",x"3397",x"0008",x"41F3", -- 07F0-07FF 
  x"46D3",x"404F",x"4000",x"A007",x"0010",x"A009",x"4377",x"003C",x"4320",x"33A0",x"0006",x"41F9",x"4377",x"33A7",x"0002",x"41F9", -- 0800-080F 
  x"0000",x"B603",x"A007",x"B501",x"2F03",x"4295",x"9002",x"B300",x"2F04",x"B501",x"2F17",x"4295",x"9009",x"B300",x"2F00",x"41FF", -- 0810-081F 
  x"0001",x"A007",x"A009",x"41FF",x"0001",x"A007",x"A00A",x"47E5",x"4287",x"B501",x"0010",x"4295",x"9FE4",x"B300",x"33AA",x"0004", -- 0820-082F 
  x"41F9",x"B501",x"4350",x"33AF",x"0001",x"41F9",x"B501",x"000F",x"A007",x"436A",x"0010",x"A007",x"B603",x"42AE",x"A00B",x"9FCC", -- 0830-083F 
  x"B200",x"4377",x"003C",x"4320",x"33B1",x"0007",x"41F9",x"42D4",x"2F00",x"A009",x"A003",x"FFA6",x"33B9",x"0005",x"4068",x"2F18", -- 0840-084F 
  x"FFFB",x"33BF",x"0008",x"478E",x"2F18",x"A00A",x"B501",x"4073",x"B501",x"4287",x"2F18",x"A009",x"A009",x"A003",x"FFF2",x"33C8", -- 0850-085F 
  x"0004",x"478E",x"B501",x"900D",x"42E7",x"B502",x"A00A",x"B502",x"A009",x"B412",x"4287",x"B412",x"4287",x"42D4",x"0001",x"428E", -- 0860-086F 
  x"8FF1",x"B300",x"B200",x"A003",x"FFEA",x"33CD",x"0004",x"478E",x"B434",x"B434",x"B501",x"9009",x"42E7",x"B603",x"A009",x"0001", -- 0870-087F 
  x"A007",x"42D4",x"0001",x"428E",x"8FF5",x"B300",x"B200",x"A003",x"FFEC",x"33D2",x"0004",x"478E",x"B412",x"B501",x"A00A",x"436A", -- 0880-088F 
  x"0001",x"A007",x"B412",x"0001",x"428E",x"B501",x"A00D",x"9FF4",x"B300",x"A003",x"FFEE",x"33D7",x"0003",x"478E",x"B603",x"429C", -- 0890-089F 
  x"9001",x"B412",x"B300",x"A003",x"FFF6",x"33DB",x"0003",x"478E",x"B603",x"42AE",x"9001",x"B412",x"B300",x"A003",x"FFF6",x"33DF", -- 08A0-08AF 
  x"0003",x"478E",x"B501",x"A00F",x"9001",x"A000",x"A003",x"FFF7",x"33E3",x"0006",x"4112",x"A017",x"A003",x"FFFA",x"33EA",x"0007", -- 08B0-08BF 
  x"4112",x"A018",x"A003",x"FFFA",x"33F2",x"0009",x"478E",x"42E7",x"A017",x"A018",x"9FFD",x"42D4",x"B300",x"A003",x"FFF5",x"33FC", -- 08C0-08CF 
  x"0001",x"4068",x"1401",x"FFFB",x"33FE",x"0001",x"4068",x"1601",x"FFFB",x"3400",x"0001",x"4068",x"1801",x"FFFB",x"3402",x"0004", -- 08D0-08DF 
  x"478E",x"0007",x"4406",x"4457",x"A009",x"444E",x"A009",x"4445",x"A009",x"443C",x"A009",x"4433",x"A009",x"442A",x"A009",x"4421", -- 08E0-08EF 
  x"A009",x"4421",x"A00A",x"443C",x"A00A",x"9001",x"A00B",x"442A",x"A00A",x"4445",x"A00A",x"A007",x"4287",x"4457",x"A00A",x"B502", -- 08F0-08FF 
  x"0000",x"4878",x"4457",x"A00A",x"B501",x"4433",x"A00A",x"442A",x"A00A",x"0000",x"B60C",x"A00A",x"B434",x"B434",x"444E",x"A00A", -- 0900-090F 
  x"4445",x"A00A",x"48C7",x"B300",x"A009",x"B300",x"B434",x"0001",x"A007",x"B434",x"0001",x"A007",x"B434",x"FFFF",x"A007",x"B501", -- 0910-091F 
  x"A00D",x"9FE7",x"B300",x"B200",x"4415",x"A003",x"FFB7",x"3407",x"0006",x"478E",x"0007",x"4406",x"4457",x"A009",x"444E",x"A009", -- 0920-092F 
  x"4445",x"A009",x"443C",x"A009",x"4433",x"A009",x"442A",x"A009",x"4421",x"A009",x"4421",x"A00A",x"442A",x"A00A",x"4445",x"A00A", -- 0930-093F 
  x"489E",x"4287",x"4457",x"A00A",x"4421",x"A00A",x"443C",x"A00A",x"4295",x"903C",x"0000",x"442A",x"A00A",x"4445",x"A00A",x"489E", -- 0940-094F 
  x"0000",x"B434",x"B502",x"B501",x"442A",x"A00A",x"429C",x"9009",x"4433",x"A00A",x"B501",x"A00A",x"B412",x"4287",x"4433",x"A009", -- 0950-095F 
  x"8001",x"0000",x"B412",x"4445",x"A00A",x"429C",x"9009",x"444E",x"A00A",x"B501",x"A00A",x"B412",x"4287",x"444E",x"A009",x"8001", -- 0960-096F 
  x"0000",x"A001",x"4457",x"A00A",x"B501",x"4287",x"4457",x"A009",x"A009",x"B434",x"B434",x"0001",x"A007",x"B603",x"428E",x"A00D", -- 0970-097F 
  x"9FD0",x"B200",x"4457",x"A00A",x"A009",x"8065",x"B412",x"0001",x"428E",x"B412",x"0001",x"442A",x"A00A",x"4445",x"A00A",x"489E", -- 0980-098F 
  x"0000",x"B434",x"B502",x"B501",x"442A",x"A00A",x"429C",x"9009",x"4433",x"A00A",x"B501",x"A00A",x"B412",x"4287",x"4433",x"A009", -- 0990-099F 
  x"8001",x"0000",x"B412",x"4445",x"A00A",x"429C",x"900A",x"444E",x"A00A",x"B501",x"A00A",x"B412",x"4287",x"444E",x"A009",x"A00B", -- 09A0-09AF 
  x"8001",x"FFFF",x"A001",x"4457",x"A00A",x"B501",x"4287",x"4457",x"A009",x"A009",x"B434",x"B434",x"0001",x"A007",x"B603",x"428E", -- 09B0-09BF 
  x"A00D",x"9FCF",x"B200",x"A00D",x"9026",x"B501",x"4457",x"A009",x"B434",x"A00B",x"B434",x"B434",x"0001",x"442A",x"A00A",x"4445", -- 09C0-09CF 
  x"A00A",x"489E",x"0000",x"B434",x"0000",x"4457",x"A00A",x"A00A",x"A00B",x"A001",x"4457",x"A00A",x"B501",x"4287",x"4457",x"A009", -- 09D0-09DF 
  x"A009",x"B434",x"B434",x"0001",x"A007",x"B603",x"428E",x"A00D",x"9FEA",x"B200",x"B300",x"4415",x"A003",x"FF39",x"340E",x"0004", -- 09E0-09EF 
  x"4112",x"A014",x"A003",x"FFFA",x"3413",x"0005",x"478E",x"0010",x"42E7",x"A014",x"42D4",x"0001",x"428E",x"B501",x"A00D",x"9FF8", -- 09F0-09FF 
  x"B200",x"A003",x"FFF1",x"3419",x"0004",x"478E",x"0000",x"B434",x"B434",x"49F7",x"A003",x"FFF7",x"341E",x"0004",x"478E",x"B502", -- 0A00-0A0F 
  x"A00F",x"9012",x"B412",x"A000",x"B412",x"B501",x"A00F",x"9006",x"A000",x"4A06",x"B412",x"A000",x"B412",x"8005",x"4A06",x"A000", -- 0A10-0A1F 
  x"B412",x"A000",x"B412",x"8008",x"B501",x"A00F",x"9004",x"A000",x"4A06",x"A000",x"8001",x"4A06",x"A003",x"FFDE",x"3423",x"0001", -- 0A20-0A2F 
  x"478E",x"4A0F",x"B412",x"B300",x"A003",x"FFF8",x"3425",x"0003",x"478E",x"4A0F",x"B300",x"A003",x"FFF9",x"3429",x"0004",x"478E", -- 0A30-0A3F 
  x"0007",x"4406",x"4457",x"A009",x"444E",x"A009",x"4445",x"A009",x"443C",x"A009",x"4433",x"A009",x"442A",x"A009",x"4421",x"A009", -- 0A40-0A4F 
  x"442A",x"A00A",x"4445",x"A00A",x"429C",x"900A",x"4421",x"A00A",x"442A",x"A00A",x"4433",x"A00A",x"0000",x"0000",x"0000",x"80E1", -- 0A50-0A5F 
  x"442A",x"A00A",x"0000",x"4433",x"A00A",x"B502",x"A007",x"A00A",x"A00B",x"B502",x"4457",x"A00A",x"A007",x"A009",x"0001",x"A007", -- 0A60-0A6F 
  x"B603",x"428E",x"A00D",x"9FEF",x"B200",x"4457",x"A00A",x"442A",x"A00A",x"A007",x"4445",x"A00A",x"428E",x"4433",x"A009",x"FFFF", -- 0A70-0A7F 
  x"4457",x"A00A",x"442A",x"A00A",x"A007",x"A009",x"0001",x"442A",x"42C9",x"442A",x"A00A",x"4445",x"A00A",x"428E",x"0000",x"4433", -- 0A80-0A8F 
  x"A00A",x"4445",x"A00A",x"A007",x"A00A",x"A00B",x"4433",x"A00A",x"4445",x"A00A",x"A007",x"0001",x"428E",x"A00A",x"A00B",x"444E", -- 0A90-0A9F 
  x"A00A",x"4445",x"A00A",x"A007",x"0001",x"428E",x"A00A",x"49F7",x"B412",x"B300",x"B501",x"4433",x"A00A",x"4445",x"A00A",x"A007", -- 0AA0-0AAF 
  x"4287",x"A009",x"0000",x"4433",x"A00A",x"444E",x"A00A",x"4445",x"A00A",x"48C7",x"B200",x"B412",x"B300",x"0000",x"4433",x"A00A", -- 0AB0-0ABF 
  x"4445",x"A00A",x"A007",x"A00A",x"A001",x"4433",x"A00A",x"4445",x"A00A",x"A007",x"A009",x"902C",x"0001",x"4445",x"A00A",x"0000", -- 0AC0-0ACF 
  x"B434",x"B502",x"4433",x"A00A",x"B502",x"A007",x"A00A",x"B412",x"444E",x"A00A",x"A007",x"A00A",x"A00B",x"A001",x"B412",x"42E7", -- 0AD0-0ADF 
  x"B502",x"4433",x"A00A",x"A007",x"A009",x"42D4",x"B434",x"B434",x"0001",x"A007",x"B603",x"428E",x"A00D",x"9FE2",x"B200",x"FFFF", -- 0AE0-0AEF 
  x"4433",x"A00A",x"4445",x"A00A",x"A007",x"4287",x"42C9",x"8FD3",x"FFFF",x"4433",x"42C9",x"0001",x"A007",x"B603",x"428E",x"A00D", -- 0AF0-0AFF 
  x"9F8E",x"B200",x"4445",x"A00A",x"0000",x"4457",x"A00A",x"B502",x"A007",x"A00A",x"A00B",x"B502",x"4457",x"A00A",x"A007",x"A009", -- 0B00-0B0F 
  x"0001",x"A007",x"B603",x"428E",x"A00D",x"9FEF",x"B200",x"4445",x"A00A",x"4457",x"A00A",x"0001",x"428E",x"A009",x"442A",x"A00A", -- 0B10-0B1F 
  x"4445",x"A00A",x"428E",x"4457",x"A00A",x"4445",x"A00A",x"A007",x"A009",x"4421",x"A00A",x"4445",x"A00A",x"4457",x"A00A",x"4421", -- 0B20-0B2F 
  x"A00A",x"443C",x"A00A",x"9001",x"A00B",x"442A",x"A00A",x"4445",x"A00A",x"428E",x"4457",x"A00A",x"4445",x"A00A",x"A007",x"0001", -- 0B30-0B3F 
  x"A007",x"4415",x"A003",x"FEF9",x"342E",x"0008",x"4068",x"2F19",x"FFFB",x"3437",x"0008",x"4068",x"2F1A",x"FFFB",x"3440",x"0008", -- 0B40-0B4F 
  x"4068",x"2F1B",x"FFFB",x"3449",x"000E",x"4068",x"2F1C",x"FFFB",x"3458",x"000C",x"4068",x"2F1D",x"FFFB",x"3465",x"0006",x"4068", -- 0B50-0B5F 
  x"2F1E",x"FFFB",x"346C",x"000D",x"478E",x"B502",x"A00D",x"9004",x"B200",x"B300",x"0000",x"8031",x"B603",x"A007",x"0001",x"428E", -- 0B60-0B6F 
  x"B501",x"A00A",x"A00D",x"A00B",x"9FF9",x"0001",x"A007",x"B502",x"489E",x"B603",x"4295",x"9004",x"B200",x"B200",x"0000",x"801D", -- 0B70-0B7F 
  x"B502",x"428E",x"B502",x"A00A",x"C000",x"A008",x"A00D",x"B502",x"0001",x"4295",x"A008",x"9003",x"B300",x"A00A",x"8009",x"B502", -- 0B80-0B8F 
  x"0001",x"428E",x"A009",x"0001",x"428E",x"404F",x"4000",x"A00E",x"B412",x"B300",x"B412",x"9001",x"A000",x"A003",x"FFC3",x"347A", -- 0B90-0B9F 
  x"000C",x"478E",x"B501",x"A00A",x"B501",x"A00F",x"9003",x"A000",x"FFFF",x"8001",x"0000",x"B434",x"B434",x"B501",x"404F",x"4000", -- 0BA0-0BAF 
  x"A008",x"9009",x"B412",x"B300",x"3FFF",x"A008",x"B501",x"A00A",x"B412",x"4287",x"8004",x"B502",x"A009",x"0001",x"B412",x"A003", -- 0BB0-0BBF 
  x"FFDE",x"3487",x"000B",x"478E",x"2F1B",x"A00A",x"B603",x"A009",x"4287",x"B603",x"A007",x"2F1B",x"A009",x"B603",x"B412",x"0000", -- 0BC0-0BCF 
  x"4878",x"B412",x"B300",x"2F1B",x"A00A",x"2F1D",x"A00A",x"429C",x"A00B",x"9002",x"0369",x"43CC",x"A003",x"FFE3",x"3493",x"0010", -- 0BD0-0BDF 
  x"478E",x"2F1A",x"A009",x"2F19",x"A009",x"2F19",x"4BA2",x"B502",x"42E7",x"2F1A",x"4BA2",x"B502",x"42D4",x"A007",x"4287",x"4BC4", -- 0BE0-0BEF 
  x"A003",x"FFEC",x"34A4",x"0002",x"478E",x"4BE1",x"492A",x"4B65",x"A003",x"FFF8",x"34A7",x"0002",x"478E",x"A000",x"4BF5",x"A003", -- 0BF0-0BFF 
  x"FFF9",x"34AA",x"0002",x"478E",x"4BE1",x"48E1",x"4B65",x"A003",x"FFF8",x"34AD",x"0007",x"4780",x"2F11",x"A00A",x"0004",x"A007", -- 0C00-0C0F 
  x"46B5",x"A003",x"FFF6",x"34B5",x"0005",x"478E",x"B501",x"A00D",x"9002",x"0000",x"43CC",x"B501",x"2F19",x"A009",x"2F19",x"4BA2", -- 0C10-0C1F 
  x"B434",x"B300",x"B502",x"A007",x"0001",x"428E",x"A00A",x"B412",x"0001",x"42AE",x"9018",x"0001",x"B502",x"A00F",x"A00B",x"9007", -- 0C20-0C2F 
  x"B412",x"B501",x"A007",x"B412",x"B501",x"4BF5",x"8FF5",x"B412",x"B300",x"B501",x"2F1E",x"A009",x"B434",x"B502",x"4C04",x"B434", -- 0C30-0C3F 
  x"B434",x"4C04",x"8004",x"B300",x"0001",x"2F1E",x"A009",x"4BE1",x"4A40",x"4B65",x"42E7",x"4B65",x"42D4",x"2F1E",x"A00A",x"0001", -- 0C40-0C4F 
  x"428E",x"9007",x"B412",x"2F1E",x"A00A",x"4C16",x"B412",x"B300",x"B412",x"A003",x"FFB8",x"34BB",x"0004",x"478E",x"0000",x"42E7", -- 0C50-0C5F 
  x"4327",x"B501",x"9007",x"4331",x"4320",x"42D4",x"B300",x"FFFF",x"42E7",x"8001",x"B300",x"4327",x"B501",x"42FE",x"A00E",x"9007", -- 0C60-0C6F 
  x"4331",x"4320",x"42D4",x"B300",x"FFFF",x"42E7",x"8001",x"B300",x"4327",x"B501",x"42FE",x"A00E",x"9003",x"4331",x"4320",x"8001", -- 0C70-0C7F 
  x"B300",x"4327",x"4331",x"4320",x"B300",x"42D4",x"B300",x"A003",x"FFD2",x"34C0",x"0002",x"478E",x"2F19",x"A009",x"2F19",x"4BA2", -- 0C80-0C8F 
  x"B434",x"9003",x"34C3",x"0001",x"41F9",x"B502",x"A007",x"0001",x"428E",x"B501",x"A00A",x"4C5E",x"B412",x"0001",x"428E",x"B412", -- 0C90-0C9F 
  x"B502",x"900A",x"0001",x"428E",x"B501",x"A00A",x"4350",x"B412",x"0001",x"428E",x"B412",x"8FF4",x"B300",x"B300",x"0020",x"4320", -- 0CA0-0CAF 
  x"A003",x"FFD7",x"34C5",x"0003",x"478E",x"B412",x"4C8C",x"4C8C",x"A003",x"FFF8",x"34C9",x"000B",x"4068",x"2F1F",x"FFFB",x"34D5", -- 0CB0-0CBF 
  x"0009",x"4068",x"2F20",x"FFFB",x"34DF",x"000D",x"478E",x"2F1B",x"A00A",x"A003",x"FFF9",x"34ED",x"000D",x"478E",x"2F1B",x"A009", -- 0CC0-0CCF 
  x"A003",x"FFF9",x"34FB",x"000B",x"478E",x"2F20",x"A00A",x"2F1F",x"A009",x"2F1B",x"A00A",x"2F20",x"A009",x"A003",x"FFF3",x"3507", -- 0CD0-0CDF 
  x"0004",x"478E",x"2F1C",x"A00A",x"2F1B",x"A009",x"4CD5",x"4CD5",x"A003",x"FFF5",x"350C",x"0003",x"478E",x"B501",x"2F19",x"A009", -- 0CE0-0CEF 
  x"2F19",x"4BA2",x"B501",x"2F19",x"428E",x"B300",x"0001",x"901A",x"B502",x"2F1B",x"A00A",x"4287",x"B412",x"4862",x"2F1B",x"A00A", -- 0CF0-0CFF 
  x"4287",x"B502",x"4287",x"2F1B",x"42C9",x"2F1B",x"A00A",x"2F1D",x"A00A",x"429C",x"A00B",x"9002",x"0369",x"43CC",x"4B65",x"B412", -- 0D00-0D0F 
  x"B300",x"8002",x"B200",x"B300",x"A003",x"FFD4",x"3510",x"0003",x"478E",x"B412",x"4CED",x"B412",x"4CED",x"A003",x"FFF7",x"3514", -- 0D10-0D1F 
  x"0002",x"478E",x"4CC7",x"B434",x"B434",x"4C16",x"B412",x"B300",x"B412",x"4CCE",x"4CED",x"A003",x"FFF2",x"3517",x"0004",x"478E", -- 0D20-0D2F 
  x"4CC7",x"B434",x"B434",x"4C16",x"B300",x"B412",x"4CCE",x"4CED",x"A003",x"FFF3",x"351C",x"0004",x"478E",x"4CC7",x"B434",x"B434", -- 0D30-0D3F 
  x"B501",x"9004",x"B412",x"B502",x"4D30",x"8FFA",x"B300",x"B412",x"4CCE",x"4CED",x"A003",x"FFEE",x"3521",x"0003",x"478E",x"4CC7", -- 0D40-0D4F 
  x"B434",x"B434",x"B603",x"4D3D",x"B434",x"B502",x"4D22",x"B434",x"B434",x"4D22",x"B434",x"4CCE",x"4D19",x"A003",x"FFED",x"3525", -- 0D50-0D5F 
  x"0007",x"478E",x"4CC7",x"B434",x"B434",x"0007",x"4406",x"442A",x"A009",x"4421",x"A009",x"0000",x"442A",x"A00A",x"9063",x"B501", -- 0D60-0D6F 
  x"4433",x"A009",x"0001",x"444E",x"A009",x"FFFF",x"4457",x"A009",x"4421",x"A00A",x"4433",x"A00A",x"A007",x"427B",x"002B",x"4295", -- 0D70-0D7F 
  x"9009",x"4433",x"A00A",x"4287",x"4433",x"A009",x"0000",x"4457",x"A009",x"8016",x"4421",x"A00A",x"4433",x"A00A",x"A007",x"427B", -- 0D80-0D8F 
  x"002D",x"4295",x"900D",x"4433",x"A00A",x"4287",x"4433",x"A009",x"0000",x"4457",x"A009",x"444E",x"A00A",x"A000",x"444E",x"A009", -- 0D90-0D9F 
  x"4457",x"A00A",x"9FD2",x"4433",x"A00A",x"442A",x"A00A",x"429C",x"9029",x"4421",x"A00A",x"4433",x"A00A",x"A007",x"427B",x"B501", -- 0DA0-0DAF 
  x"9015",x"454C",x"A00B",x"9007",x"B300",x"442A",x"A00A",x"A000",x"442A",x"A009",x"800A",x"B412",x"2F08",x"A00A",x"4C04",x"4BF5", -- 0DB0-0DBF 
  x"4433",x"A00A",x"4287",x"4433",x"A009",x"8005",x"B300",x"4433",x"A00A",x"442A",x"A009",x"4433",x"A00A",x"442A",x"A00A",x"429C", -- 0DC0-0DCF 
  x"A00B",x"9FD7",x"444E",x"A00A",x"A00F",x"9001",x"A000",x"4433",x"A00A",x"442A",x"A00A",x"428E",x"B501",x"9006",x"B300",x"4421", -- 0DD0-0DDF 
  x"A00A",x"4433",x"A00A",x"A007",x"4415",x"B434",x"4CCE",x"B412",x"4CED",x"B412",x"A003",x"FF73",x"352D",x"0002",x"0022",x"41D8", -- 0DE0-0DEF 
  x"4D62",x"B300",x"A003",x"FFF8",x"3530",x"0002",x"478E",x"4CC7",x"B434",x"B434",x"0004",x"4406",x"B501",x"A00F",x"9002",x"0012", -- 0DF0-0DFF 
  x"43CC",x"0002",x"443C",x"A009",x"4433",x"A009",x"442A",x"A009",x"0001",x"4433",x"A00A",x"443C",x"A00A",x"4A0F",x"4433",x"A009", -- 0E00-0E0F 
  x"9003",x"442A",x"A00A",x"4C04",x"4433",x"A00A",x"9008",x"442A",x"A00A",x"442A",x"A00A",x"4C04",x"442A",x"A009",x"8FEA",x"4415", -- 0E10-0E1F 
  x"B412",x"4CCE",x"4CED",x"A003",x"FFCF",x"3533",x"0002",x"478E",x"2F08",x"A00A",x"0010",x"4295",x"9002",x"4C8C",x"802C",x"4CC7", -- 0E20-0E2F 
  x"B412",x"B501",x"A00F",x"9004",x"A000",x"3536",x"0001",x"41F9",x"B501",x"A00D",x"9005",x"3538",x"0002",x"41F9",x"B300",x"801A", -- 0E30-0E3F 
  x"FFFF",x"B412",x"B501",x"9004",x"2F08",x"A00A",x"4C16",x"8FFA",x"B300",x"B501",x"A00F",x"A00B",x"900A",x"0030",x"A007",x"B501", -- 0E40-0E4F 
  x"0039",x"42AE",x"9002",x"0007",x"A007",x"4320",x"8FF2",x"0020",x"4320",x"B300",x"4CCE",x"A003",x"FFC8",x"353B",x"0003",x"478E", -- 0E50-0E5F 
  x"B412",x"4E28",x"4E28",x"A003",x"FFF8",x"353F",x"0006",x"478E",x"3FFF",x"A008",x"B501",x"4287",x"B412",x"A00A",x"A003",x"FFF5", -- 0E60-0E6F 
  x"3546",x"0004",x"478E",x"48B2",x"B501",x"404F",x"4000",x"429C",x"9003",x"B300",x"0000",x"800A",x"4E68",x"B412",x"B300",x"404F", -- 0E70-0E7F 
  x"4000",x"429C",x"9002",x"0000",x"8001",x"FFFF",x"A003",x"FFE8",x"354B",x"0001",x"478E",x"B502",x"4E73",x"9011",x"B412",x"4E68", -- 0E80-0E8F 
  x"3FFF",x"A008",x"B434",x"B603",x"42AE",x"9005",x"B412",x"B300",x"A007",x"A00A",x"8003",x"B200",x"B300",x"0000",x"8003",x"9002", -- 0E90-0E9F 
  x"B300",x"0000",x"A003",x"FFE4",x"354D",x"0001",x"478E",x"B603",x"4E8B",x"A003",x"FFF9",x"354F",x"0001",x"478E",x"B501",x"42E7", -- 0EA0-0EAF 
  x"B434",x"B434",x"B502",x"4E73",x"A00D",x"B502",x"A00D",x"A008",x"42D4",x"4E73",x"A00D",x"A008",x"9002",x"B200",x"806F",x"B502", -- 0EB0-0EBF 
  x"4E73",x"A00D",x"9017",x"B501",x"4287",x"4BC4",x"B434",x"B502",x"A009",x"404F",x"4000",x"B502",x"0001",x"428E",x"42C9",x"B501", -- 0EC0-0ECF 
  x"42E7",x"A007",x"A009",x"42D4",x"0001",x"428E",x"404F",x"4000",x"A007",x"8054",x"B502",x"4E68",x"3FFF",x"A008",x"B434",x"B603", -- 0ED0-0EDF 
  x"42AE",x"9008",x"B412",x"B300",x"B434",x"42E7",x"A007",x"A009",x"42D4",x"801B",x"B501",x"4287",x"4BC4",x"B412",x"42E7",x"B501", -- 0EE0-0EEF 
  x"42E7",x"B412",x"4862",x"B300",x"42D4",x"404F",x"4000",x"B502",x"0001",x"428E",x"42C9",x"B412",x"B502",x"42D4",x"A007",x"A009", -- 0EF0-0EFF 
  x"0001",x"428E",x"404F",x"4000",x"A007",x"4E68",x"3FFF",x"A008",x"B603",x"A007",x"0001",x"428E",x"A00A",x"A00D",x"B502",x"0001", -- 0F00-0F0F 
  x"42AE",x"A008",x"9003",x"0001",x"428E",x"8FF2",x"B502",x"A00A",x"4E73",x"A00D",x"B502",x"0001",x"4295",x"A008",x"9003",x"B300", -- 0F10-0F1F 
  x"A00A",x"800C",x"B412",x"0001",x"428E",x"B412",x"404F",x"4000",x"A007",x"B502",x"A009",x"404F",x"4000",x"A007",x"A003",x"FF7B", -- 0F20-0F2F 
  x"3551",x"0002",x"478E",x"B501",x"4E73",x"9017",x"3554",x"0002",x"41F9",x"4E68",x"3FFF",x"A008",x"B502",x"A007",x"B412",x"B603", -- 0F30-0F3F 
  x"42AE",x"9006",x"B501",x"A00A",x"4F33",x"0001",x"A007",x"8FF7",x"B200",x"3557",x"0002",x"41F9",x"8001",x"4E28",x"A003",x"FFE0", -- 0F40-0F4F 
  x"355A",x"0006",x"4068",x"2F21",x"FFFB",x"3561",x"0001",x"478E",x"2F21",x"A00A",x"2801",x"A00A",x"2F21",x"A009",x"A003",x"FFF5", -- 0F50-0F5F 
  x"3563",x"0001",x"478E",x"0000",x"2801",x"A00A",x"0001",x"428E",x"2F21",x"A00A",x"428E",x"900A",x"2801",x"A00A",x"0002",x"428E", -- 0F60-0F6F 
  x"2F21",x"A00A",x"428E",x"B434",x"4EAE",x"8FEE",x"B412",x"2F21",x"A009",x"A003",x"FFE5",x"3565",x"0005",x"478E",x"B501",x"4E73", -- 0F70-0F7F 
  x"901C",x"B501",x"42E7",x"4E68",x"3FFF",x"A008",x"B412",x"B502",x"A007",x"FFFF",x"A007",x"B412",x"B501",x"900C",x"B412",x"B501", -- 0F80-0F8F 
  x"A00A",x"4F7E",x"B502",x"A009",x"FFFF",x"A007",x"B412",x"FFFF",x"A007",x"8FF2",x"B200",x"42D4",x"8001",x"4CED",x"A003",x"FFDB", -- 0F90-0F9F 
  x"356B",x"0007",x"478E",x"B501",x"4E73",x"902A",x"4E68",x"3FFF",x"A008",x"B501",x"9023",x"B412",x"4377",x"B502",x"436A",x"B501", -- 0FA0-0FAF 
  x"436A",x"B501",x"A00A",x"B501",x"436A",x"B501",x"48B2",x"404F",x"4000",x"429C",x"9005",x"FFFF",x"436A",x"FFFF",x"436A",x"8005", -- 0FB0-0FBF 
  x"B501",x"48B2",x"4E68",x"436A",x"436A",x"B501",x"4F33",x"4FA3",x"0001",x"A007",x"B412",x"FFFF",x"A007",x"8FDB",x"B200",x"8001", -- 0FC0-0FCF 
  x"B300",x"A003",x"FFCD",x"3573",x"000B",x"478E",x"0008",x"4406",x"4CC7",x"4421",x"A009",x"442A",x"A009",x"0001",x"442A",x"A00A", -- 0FD0-0FDF 
  x"4433",x"A009",x"FFFF",x"4433",x"42C9",x"4460",x"A009",x"0000",x"444E",x"A009",x"0000",x"4457",x"A009",x"B501",x"4433",x"A00A", -- 0FE0-0FEF 
  x"4E8B",x"4433",x"A00A",x"4E8B",x"442A",x"A00A",x"443C",x"A009",x"FFFF",x"443C",x"42C9",x"B502",x"443C",x"A00A",x"4E8B",x"4433", -- 0FF0-0FFF 
  x"A00A",x"4E8B",x"444E",x"A00A",x"443C",x"A00A",x"B434",x"4EAE",x"444E",x"A009",x"B502",x"4433",x"A00A",x"4E8B",x"443C",x"A00A", -- 1000-100F 
  x"4E8B",x"4457",x"A00A",x"443C",x"A00A",x"B434",x"4EAE",x"4457",x"A009",x"443C",x"A00A",x"A00D",x"9FDB",x"444E",x"A00A",x"4433", -- 1010-101F 
  x"A00A",x"4E8B",x"4460",x"A00A",x"4BF5",x"444E",x"A00A",x"4433",x"A00A",x"B434",x"4EAE",x"444E",x"A009",x"4457",x"A00A",x"4433", -- 1020-102F 
  x"A00A",x"4E8B",x"4460",x"A00A",x"4BFD",x"4457",x"A00A",x"4433",x"A00A",x"B434",x"4EAE",x"4457",x"A009",x"442A",x"A00A",x"443C", -- 1030-103F 
  x"A009",x"FFFF",x"443C",x"42C9",x"B502",x"443C",x"A00A",x"4E8B",x"442A",x"A00A",x"4445",x"A009",x"FFFF",x"4445",x"42C9",x"4CC7", -- 1040-104F 
  x"B434",x"B434",x"B412",x"B502",x"4445",x"A00A",x"4E8B",x"B502",x"4C04",x"444E",x"A00A",x"443C",x"A00A",x"4E8B",x"4457",x"A00A", -- 1050-105F 
  x"4445",x"A00A",x"4E8B",x"4C04",x"4BFD",x"4460",x"A00A",x"4D22",x"B43C",x"B412",x"4CCE",x"B412",x"4CED",x"B412",x"4445",x"A00A", -- 1060-106F 
  x"B434",x"4EAE",x"4445",x"A00A",x"A00D",x"9FD6",x"B434",x"443C",x"A00A",x"B434",x"4EAE",x"B412",x"443C",x"A00A",x"A00D",x"9FC1", -- 1070-107F 
  x"4CED",x"4421",x"A00A",x"4CCE",x"B412",x"4F7E",x"B412",x"4CED",x"4433",x"A00A",x"A00D",x"9F56",x"4415",x"A003",x"FF44",x"357F", -- 1080-108F 
  x"0011",x"478E",x"0003",x"4406",x"4421",x"A009",x"0000",x"4421",x"A00A",x"442A",x"A009",x"442A",x"A00A",x"B501",x"9023",x"0001", -- 1090-109F 
  x"428E",x"442A",x"A009",x"442A",x"A00A",x"4EA7",x"4421",x"A00A",x"4433",x"A009",x"4433",x"A00A",x"B501",x"9011",x"0001",x"428E", -- 10A0-10AF 
  x"4433",x"A009",x"4433",x"A00A",x"442A",x"A00A",x"0001",x"A007",x"4433",x"A00A",x"0001",x"A007",x"4DF7",x"4EAE",x"8FEB",x"B300", -- 10B0-10BF 
  x"4EAE",x"8FD9",x"B300",x"4415",x"A003",x"FFC9",x"3591",x"0005",x"478E",x"2F11",x"A00A",x"B501",x"4287",x"A00A",x"B502",x"0002", -- 10C0-10CF 
  x"A007",x"A00A",x"433F",x"0020",x"4320",x"B501",x"A00A",x"9004",x"B501",x"A00A",x"A007",x"8FEF",x"B300",x"A003",x"FFE7",x"3597", -- 10D0-10DF 
  x"0005",x"478E",x"2F11",x"A00A",x"B501",x"436A",x"B501",x"4287",x"A00A",x"B502",x"0002",x"A007",x"A00A",x"433F",x"0020",x"4320", -- 10E0-10EF 
  x"B501",x"A00A",x"9004",x"B501",x"A00A",x"A007",x"8FED",x"B300",x"A003",x"FFE5",x"359D",x"0006",x"4068",x"A003",x"FFFB",x"35A4", -- 10F0-10FF 
  x"0008",x"478E",x"43F0",x"0020",x"45F2",x"466C",x"B501",x"9012",x"46AC",x"B300",x"4287",x"41FF",x"B412",x"2F0F",x"A009",x"B501", -- 1100-110F 
  x"46B5",x"404F",x"A003",x"4307",x"2F0F",x"A009",x"0001",x"2F10",x"A009",x"8003",x"B200",x"0003",x"43CC",x"A003",x"FFE0",x"35AD", -- 1110-111F 
  x"0006",x"478E",x"0020",x"45F2",x"466C",x"900E",x"2F0F",x"A009",x"41FF",x"B501",x"A00A",x"A007",x"2F11",x"A009",x"41FF",x"4287", -- 1120-112F 
  x"A00A",x"2F13",x"A009",x"8004",x"B300",x"35B4",x"000F",x"41F9",x"A003",x"FFE5",x"35C4",x"000A",x"478E",x"4377",x"B501",x"0000", -- 1130-113F 
  x"4295",x"9003",x"35CF",x"0013",x"41F9",x"B501",x"0003",x"4295",x"9003",x"35E3",x"0014",x"41F9",x"B501",x"0006",x"4295",x"9003", -- 1140-114F 
  x"35F8",x"0014",x"41F9",x"B501",x"0009",x"4295",x"9003",x"360D",x"0030",x"41F9",x"B501",x"0012",x"4295",x"9003",x"363E",x"0012", -- 1150-115F 
  x"41F9",x"B501",x"0369",x"4295",x"9003",x"3651",x"0013",x"41F9",x"B501",x"1234",x"4295",x"9003",x"3665",x"004C",x"41F9",x"A003", -- 1160-116F 
  x"FFC9",x"36B2",x"0005",x"478E",x"47AE",x"41FF",x"0003",x"428E",x"B501",x"436A",x"A00A",x"4287",x"B501",x"436A",x"A00A",x"B501", -- 1170-117F 
  x"436A",x"0040",x"428E",x"41FF",x"B412",x"0007",x"A008",x"0018",x"A007",x"A009",x"A003",x"FFE5",x"36B8",x"0002",x"478E",x"0007", -- 1180-118F 
  x"4320",x"36BB",x"0008",x"41F9",x"A003",x"FFF6",x"36C4",x"0002",x"478E",x"0007",x"4320",x"36C7",x"0004",x"41F9",x"4720",x"A003", -- 1190-119F 
  x"FFF5",x"36CC",x"0002",x"478E",x"36CF",x"0029",x"41F9",x"4377",x"FA00",x"0100",x"44E0",x"46D3",x"36F9",x"0002",x"41F9",x"A003", -- 11A0-11AF 
  x"FFF0",x"36FC",x"0005",x"478E",x"2F09",x"A00A",x"0100",x"44E0",x"A003",x"FFF7",x"3702",x"0007",x"4780",x"003C",x"4320",x"370A", -- 11B0-11BF 
  x"0004",x"41F9",x"4377",x"51B4",x"370F",x"0007",x"41F3",x"4638",x"9FF9",x"003C",x"4320",x"3717",x"0003",x"41F9",x"A003",x"FFEA", -- 11C0-11CF 
  x"371B",x"0003",x"478E",x"0010",x"2F08",x"A009",x"A003",x"FFF8",x"371F",x"0007",x"478E",x"000A",x"2F08",x"A009",x"A003",x"FFF8", -- 11D0-11DF 
  x"3727",x"0005",x"478E",x"B501",x"3FFF",x"42AE",x"B502",x"C000",x"429C",x"A00E",x"9002",x"1234",x"43CC",x"4307",x"A003",x"51E3", -- 11E0-11EF 
  x"A003",x"4D62",x"A003",x"FFEC",x"372D",x"0002",x"478E",x"436A",x"A003",x"FFFA",x"3730",x"0002",x"478E",x"A007",x"A003",x"FFFA", -- 11F0-11FF 
  x"3733",x"0002",x"478E",x"428E",x"A003",x"FFFA",x"3736",x"0002",x"478E",x"42B5",x"A003",x"FFFA",x"3739",x"0002",x"478E",x"4A31", -- 1200-120F 
  x"A003",x"FFFA",x"373C",x"0005",x"478E",x"4A0F",x"A003",x"FFFA",x"3742",x"0004",x"478E",x"4A39",x"A003",x"FFFA",x"3747",x"0001", -- 1210-121F 
  x"478E",x"4F33",x"A003",x"FFFA",x"3749",x"0001",x"478E",x"4BF5",x"A003",x"FFFA",x"374B",x"0001",x"478E",x"4BFD",x"A003",x"FFFA", -- 1220-122F 
  x"374D",x"0001",x"478E",x"4C04",x"A003",x"FFFA",x"374F",x"0001",x"478E",x"4D22",x"A003",x"FFFA",x"3751",x"0004",x"478E",x"4C16", -- 1230-123F 
  x"47AE",x"47AE",x"4A39",x"4D30",x"A003",x"FFF6",x"3756",x"0003",x"478E",x"4D3D",x"A003",x"FFFA",x"375A",x"0002",x"478E",x"4D4F", -- 1240-124F 
  x"A003",x"FFFA",x"375D",x"0001",x"478E",x"4DF7",x"A003",x"FFFA",x"375F",x"0001",x"478E",x"A00A",x"5221",x"A003",x"0000",x"2F00", -- 1250-125F 
  SHA(10*16-1 downto 9*16),
  SHA(9*16-1 downto 8*16),
  SHA(8*16-1 downto 7*16),
  SHA(7*16-1 downto 6*16),
  SHA(6*16-1 downto 5*16),
  SHA(5*16-1 downto 4*16),
  SHA(4*16-1 downto 3*16),
  SHA(3*16-1 downto 2*16),
  SHA(2*16-1 downto 1*16),
  SHA(1*16-1 downto 0*16),
  others=>x"0000");

-- Textspeicher
type ByteRAMTYPE is array(0 to 4*1024-1) of STD_LOGIC_VECTOR (7 downto 0);
signal ByteRAM: ByteRAMTYPE:=(
  x"28",x"20",x"7B",x"20",x"7D",x"20",x"43",x"4F",x"4D",x"50",x"49",x"4C",x"45",x"20",x"28",x"4C", -- 3000-300F 
  x"49",x"54",x"2C",x"29",x"20",x"4C",x"49",x"54",x"2C",x"20",x"28",x"43",x"4F",x"4E",x"53",x"54", -- 3010-301F 
  x"41",x"4E",x"54",x"3A",x"29",x"20",x"43",x"4F",x"4E",x"53",x"54",x"41",x"4E",x"54",x"20",x"4B", -- 3020-302F 
  x"45",x"59",x"41",x"44",x"52",x"20",x"53",x"50",x"20",x"52",x"50",x"20",x"50",x"43",x"20",x"58", -- 3030-303F 
  x"42",x"49",x"54",x"20",x"53",x"4D",x"55",x"44",x"47",x"45",x"42",x"49",x"54",x"20",x"52",x"50", -- 3040-304F 
  x"30",x"20",x"49",x"52",x"41",x"4D",x"41",x"44",x"52",x"20",x"4A",x"52",x"41",x"4D",x"41",x"44", -- 3050-305F 
  x"52",x"20",x"58",x"4F",x"46",x"46",x"20",x"43",x"52",x"42",x"5A",x"45",x"49",x"47",x"20",x"43", -- 3060-306F 
  x"52",x"44",x"50",x"20",x"42",x"41",x"53",x"45",x"20",x"54",x"49",x"42",x"20",x"49",x"4E",x"31", -- 3070-307F 
  x"20",x"49",x"4E",x"32",x"20",x"49",x"4E",x"33",x"20",x"49",x"4E",x"34",x"20",x"45",x"52",x"52", -- 3080-308F 
  x"4F",x"52",x"4E",x"52",x"20",x"44",x"50",x"20",x"53",x"54",x"41",x"54",x"20",x"4C",x"46",x"41", -- 3090-309F 
  x"20",x"42",x"41",x"4E",x"46",x"20",x"42",x"5A",x"45",x"49",x"47",x"20",x"44",x"50",x"4D",x"45", -- 30A0-30AF 
  x"52",x"4B",x"20",x"43",x"53",x"50",x"20",x"4C",x"4F",x"43",x"41",x"4C",x"41",x"44",x"44",x"52", -- 30B0-30BF 
  x"20",x"4C",x"4F",x"43",x"41",x"4C",x"41",x"44",x"52",x"45",x"53",x"53",x"45",x"20",x"56",x"45", -- 30C0-30CF 
  x"52",x"53",x"49",x"4F",x"4E",x"20",x"52",x"45",x"54",x"55",x"52",x"4E",x"20",x"28",x"4D",x"43", -- 30D0-30DF 
  x"4F",x"44",x"45",x"3A",x"29",x"20",x"4D",x"43",x"4F",x"44",x"45",x"20",x"4D",x"49",x"4E",x"55", -- 30E0-30EF 
  x"53",x"20",x"55",x"2B",x"20",x"55",x"2A",x"20",x"30",x"3D",x"20",x"30",x"4C",x"54",x"20",x"45", -- 30F0-30FF 
  x"4D",x"49",x"54",x"43",x"4F",x"44",x"45",x"20",x"4E",x"4F",x"54",x"20",x"41",x"4E",x"44",x"20", -- 3100-310F 
  x"4F",x"52",x"20",x"4B",x"45",x"59",x"43",x"4F",x"44",x"45",x"20",x"2B",x"20",x"21",x"20",x"40", -- 3110-311F 
  x"20",x"53",x"57",x"41",x"50",x"20",x"4F",x"56",x"45",x"52",x"20",x"44",x"55",x"50",x"20",x"52", -- 3120-312F 
  x"4F",x"54",x"20",x"44",x"52",x"4F",x"50",x"20",x"32",x"53",x"57",x"41",x"50",x"20",x"32",x"4F", -- 3130-313F 
  x"56",x"45",x"52",x"20",x"32",x"44",x"55",x"50",x"20",x"32",x"44",x"52",x"4F",x"50",x"20",x"4E", -- 3140-314F 
  x"4F",x"4F",x"50",x"20",x"42",x"2C",x"20",x"5A",x"2C",x"20",x"28",x"57",x"4F",x"52",x"44",x"3A", -- 3150-315F 
  x"29",x"20",x"57",x"4F",x"52",x"44",x"3A",x"20",x"22",x"20",x"2E",x"22",x"20",x"48",x"45",x"52", -- 3160-316F 
  x"45",x"20",x"4A",x"52",x"42",x"49",x"54",x"20",x"4A",x"52",x"30",x"42",x"49",x"54",x"20",x"58", -- 3170-317F 
  x"53",x"45",x"54",x"42",x"54",x"20",x"41",x"4C",x"4C",x"4F",x"54",x"20",x"42",x"52",x"41",x"4E", -- 3180-318F 
  x"43",x"48",x"2C",x"20",x"30",x"42",x"52",x"41",x"4E",x"43",x"48",x"2C",x"20",x"42",x"45",x"47", -- 3190-319F 
  x"49",x"4E",x"20",x"41",x"47",x"41",x"49",x"4E",x"20",x"55",x"4E",x"54",x"49",x"4C",x"20",x"49", -- 31A0-31AF 
  x"46",x"20",x"45",x"4E",x"44",x"5F",x"49",x"46",x"20",x"45",x"4C",x"53",x"45",x"20",x"57",x"48", -- 31B0-31BF 
  x"49",x"4C",x"45",x"20",x"52",x"45",x"50",x"45",x"41",x"54",x"20",x"43",x"40",x"20",x"43",x"21", -- 31C0-31CF 
  x"20",x"31",x"2B",x"20",x"2D",x"20",x"3D",x"20",x"4C",x"54",x"20",x"3E",x"20",x"2A",x"20",x"42", -- 31D0-31DF 
  x"59",x"45",x"20",x"42",x"59",x"45",x"20",x"20",x"2B",x"21",x"20",x"52",x"3E",x"20",x"3E",x"52", -- 31E0-31EF 
  x"20",x"52",x"20",x"2C",x"20",x"45",x"58",x"45",x"43",x"55",x"54",x"45",x"20",x"4B",x"45",x"59", -- 31F0-31FF 
  x"20",x"45",x"4D",x"49",x"54",x"20",x"53",x"48",x"4C",x"31",x"36",x"20",x"44",x"49",x"47",x"20", -- 3200-320F 
  x"54",x"59",x"50",x"45",x"20",x"48",x"47",x"2E",x"20",x"48",x"2E",x"20",x"2E",x"20",x"3F",x"20", -- 3210-321F 
  x"43",x"52",x"20",x"66",x"6C",x"3E",x"20",x"2F",x"66",x"6C",x"3E",x"20",x"66",x"72",x"3E",x"20", -- 3220-322F 
  x"2F",x"66",x"72",x"3E",x"20",x"46",x"45",x"48",x"4C",x"45",x"52",x"54",x"45",x"58",x"54",x"20", -- 3230-323F 
  x"44",x"49",x"53",x"41",x"42",x"4C",x"45",x"20",x"77",x"65",x"69",x"74",x"65",x"72",x"20",x"6E", -- 3240-324F 
  x"61",x"63",x"68",x"20",x"54",x"61",x"73",x"74",x"65",x"20",x"45",x"53",x"43",x"41",x"50",x"45", -- 3250-325F 
  x"20",x"20",x"45",x"52",x"52",x"4F",x"52",x"20",x"3F",x"3F",x"3F",x"20",x"46",x"45",x"48",x"4C", -- 3260-326F 
  x"45",x"52",x"54",x"45",x"58",x"54",x"20",x"45",x"52",x"52",x"4F",x"52",x"20",x"2D",x"20",x"46", -- 3270-327F 
  x"65",x"68",x"6C",x"65",x"72",x"20",x"4E",x"75",x"6D",x"6D",x"65",x"72",x"20",x"20",x"43",x"53", -- 3280-328F 
  x"50",x"21",x"20",x"43",x"53",x"50",x"3F",x"20",x"4C",x"4F",x"43",x"41",x"4C",x"20",x"45",x"4E", -- 3290-329F 
  x"44",x"5F",x"4C",x"4F",x"43",x"41",x"4C",x"20",x"4C",x"30",x"20",x"4C",x"31",x"20",x"4C",x"32", -- 32A0-32AF 
  x"20",x"4C",x"33",x"20",x"4C",x"34",x"20",x"4C",x"35",x"20",x"4C",x"36",x"20",x"4C",x"37",x"20", -- 32B0-32BF 
  x"27",x"20",x"49",x"4E",x"43",x"52",x"34",x"20",x"4B",x"45",x"59",x"5F",x"49",x"4E",x"54",x"20", -- 32C0-32CF 
  x"4B",x"45",x"59",x"43",x"4F",x"44",x"45",x"32",x"20",x"45",x"58",x"50",x"45",x"43",x"54",x"20", -- 32D0-32DF 
  x"44",x"49",x"47",x"49",x"54",x"20",x"4E",x"55",x"4D",x"42",x"45",x"52",x"20",x"57",x"4F",x"52", -- 32E0-32EF 
  x"44",x"20",x"5A",x"3D",x"20",x"46",x"49",x"4E",x"44",x"20",x"4C",x"43",x"46",x"41",x"20",x"43", -- 32F0-32FF 
  x"4F",x"4D",x"50",x"49",x"4C",x"45",x"2C",x"20",x"43",x"52",x"45",x"41",x"54",x"45",x"20",x"49", -- 3300-330F 
  x"4E",x"54",x"45",x"52",x"50",x"52",x"45",x"54",x"20",x"51",x"55",x"49",x"54",x"20",x"2F",x"6F", -- 3310-331F 
  x"6B",x"3E",x"20",x"6F",x"6B",x"20",x"6F",x"6B",x"3E",x"20",x"2F",x"6F",x"6B",x"3E",x"20",x"6F", -- 3320-332F 
  x"6B",x"20",x"53",x"54",x"41",x"52",x"54",x"20",x"46",x"4F",x"52",x"54",x"59",x"2D",x"46",x"4F", -- 3330-333F 
  x"52",x"54",x"48",x"20",x"53",x"4D",x"55",x"44",x"47",x"45",x"20",x"28",x"49",x"4D",x"4D",x"45", -- 3340-334F 
  x"44",x"49",x"41",x"54",x"45",x"3A",x"29",x"20",x"28",x"43",x"4F",x"4D",x"50",x"49",x"4C",x"45", -- 3350-335F 
  x"3A",x"29",x"20",x"28",x"3A",x"29",x"20",x"49",x"4D",x"4D",x"45",x"44",x"49",x"41",x"54",x"45", -- 3360-336F 
  x"3A",x"20",x"43",x"4F",x"4D",x"50",x"49",x"4C",x"45",x"3A",x"20",x"3A",x"20",x"3B",x"20",x"44", -- 3370-337F 
  x"55",x"42",x"49",x"54",x"20",x"4C",x"47",x"2E",x"20",x"4E",x"47",x"2E",x"20",x"78",x"20",x"2C", -- 3380-338F 
  x"20",x"44",x"55",x"4D",x"50",x"5A",x"20",x"27",x"20",x"53",x"54",x"41",x"52",x"54",x"20",x"20", -- 3390-339F 
  x"44",x"55",x"4D",x"50",x"5A",x"3E",x"20",x"20",x"20",x"20",x"20",x"2D",x"2D",x"20",x"20",x"2D", -- 33A0-33AF 
  x"20",x"2F",x"44",x"55",x"4D",x"50",x"5A",x"3E",x"20",x"52",x"41",x"4D",x"50",x"31",x"20",x"56", -- 33B0-33BF 
  x"41",x"52",x"49",x"41",x"42",x"4C",x"45",x"20",x"4D",x"4F",x"56",x"45",x"20",x"46",x"49",x"4C", -- 33C0-33CF 
  x"4C",x"20",x"44",x"55",x"4D",x"50",x"20",x"4D",x"41",x"58",x"20",x"4D",x"49",x"4E",x"20",x"41", -- 33D0-33DF 
  x"42",x"53",x"20",x"4D",x"55",x"4C",x"54",x"5F",x"49",x"20",x"4D",x"55",x"4C",x"54",x"5F",x"49", -- 33E0-33EF 
  x"49",x"20",x"53",x"55",x"50",x"45",x"52",x"4D",x"55",x"4C",x"54",x"20",x"41",x"20",x"42",x"20", -- 33F0-33FF 
  x"43",x"20",x"53",x"4D",x"55",x"4C",x"20",x"41",x"44",x"44",x"49",x"45",x"52",x"20",x"44",x"49", -- 3400-340F 
  x"33",x"32",x"20",x"44",x"49",x"56",x"33",x"32",x"20",x"2F",x"4D",x"4F",x"44",x"20",x"2F",x"4D", -- 3410-341F 
  x"4F",x"44",x"20",x"2F",x"20",x"4D",x"4F",x"44",x"20",x"53",x"44",x"49",x"56",x"20",x"4F",x"50", -- 3420-342F 
  x"45",x"52",x"41",x"4E",x"44",x"31",x"20",x"4F",x"50",x"45",x"52",x"41",x"4E",x"44",x"32",x"20", -- 3430-343F 
  x"45",x"52",x"47",x"45",x"42",x"4E",x"49",x"53",x"20",x"5A",x"41",x"48",x"4C",x"45",x"4E",x"53", -- 3440-344F 
  x"50",x"45",x"49",x"43",x"48",x"45",x"52",x"20",x"53",x"50",x"45",x"49",x"43",x"48",x"45",x"52", -- 3450-345F 
  x"45",x"4E",x"44",x"45",x"20",x"53",x"43",x"48",x"49",x"45",x"42",x"20",x"53",x"4C",x"58",x"2D", -- 3460-346F 
  x"3E",x"45",x"52",x"47",x"45",x"42",x"4E",x"49",x"53",x"20",x"4F",x"50",x"45",x"52",x"41",x"4E", -- 3470-347F 
  x"44",x"2D",x"3E",x"53",x"4C",x"58",x"20",x"53",x"50",x"45",x"49",x"43",x"48",x"45",x"52",x"48", -- 3480-348F 
  x"4F",x"4C",x"20",x"32",x"4F",x"50",x"45",x"52",x"41",x"4E",x"44",x"45",x"4E",x"2D",x"3E",x"32", -- 3490-349F 
  x"53",x"4C",x"58",x"20",x"4E",x"2B",x"20",x"4E",x"2D",x"20",x"4E",x"2A",x"20",x"52",x"45",x"43", -- 34A0-34AF 
  x"55",x"52",x"53",x"45",x"20",x"4E",x"2F",x"4D",x"4F",x"44",x"20",x"48",x"47",x"30",x"2E",x"20", -- 34B0-34BF 
  x"4E",x"2E",x"20",x"2D",x"20",x"4E",x"42",x"2E",x"20",x"42",x"4C",x"4F",x"43",x"4B",x"41",x"4E", -- 34C0-34CF 
  x"46",x"41",x"4E",x"47",x"20",x"42",x"4C",x"4F",x"43",x"4B",x"45",x"4E",x"44",x"45",x"20",x"4E", -- 34D0-34DF 
  x"45",x"42",x"45",x"4E",x"52",x"45",x"43",x"48",x"4E",x"55",x"4E",x"47",x"20",x"48",x"41",x"55", -- 34E0-34EF 
  x"50",x"54",x"52",x"45",x"43",x"48",x"4E",x"55",x"4E",x"47",x"20",x"52",x"45",x"43",x"48",x"45", -- 34F0-34FF 
  x"4E",x"42",x"4C",x"4F",x"43",x"4B",x"20",x"49",x"4E",x"49",x"54",x"20",x"41",x"2B",x"30",x"20", -- 3500-350F 
  x"42",x"2B",x"30",x"20",x"4E",x"2F",x"20",x"4E",x"4D",x"4F",x"44",x"20",x"4E",x"47",x"47",x"54", -- 3510-351F 
  x"20",x"4E",x"42",x"4B",x"20",x"4E",x"4E",x"55",x"4D",x"42",x"45",x"52",x"20",x"4E",x"22",x"20", -- 3520-352F 
  x"4E",x"5E",x"20",x"4E",x"2E",x"20",x"2D",x"20",x"30",x"20",x"20",x"4E",x"42",x"2E",x"20",x"5A", -- 3530-353F 
  x"45",x"52",x"4C",x"45",x"47",x"20",x"4F",x"42",x"4A",x"3F",x"20",x"4C",x"20",x"47",x"20",x"48", -- 3540-354F 
  x"20",x"4F",x"2E",x"20",x"5B",x"20",x"20",x"5D",x"20",x"20",x"53",x"50",x"4D",x"45",x"52",x"4B", -- 3550-355F 
  x"20",x"5B",x"20",x"5D",x"20",x"4F",x"42",x"4A",x"2B",x"30",x"20",x"4F",x"42",x"4A",x"44",x"55", -- 3560-356F 
  x"4D",x"50",x"20",x"49",x"4E",x"56",x"45",x"52",x"54",x"49",x"45",x"52",x"45",x"4E",x"20",x"56", -- 3570-357F 
  x"41",x"4E",x"44",x"45",x"52",x"4D",x"4F",x"4E",x"44",x"45",x"4D",x"41",x"54",x"52",x"49",x"58", -- 3580-358F 
  x"20",x"56",x"4C",x"49",x"53",x"54",x"20",x"57",x"4C",x"49",x"53",x"54",x"20",x"52",x"45",x"54", -- 3590-359F 
  x"55",x"52",x"4E",x"20",x"52",x"45",x"50",x"4C",x"41",x"43",x"45",x"3A",x"20",x"46",x"4F",x"52", -- 35A0-35AF 
  x"47",x"45",x"54",x"20",x"6E",x"69",x"63",x"68",x"74",x"20",x"67",x"65",x"66",x"75",x"6E",x"64", -- 35B0-35BF 
  x"65",x"6E",x"20",x"20",x"46",x"45",x"48",x"4C",x"45",x"52",x"54",x"45",x"58",x"54",x"20",x"44", -- 35C0-35CF 
  x"69",x"76",x"69",x"73",x"69",x"6F",x"6E",x"20",x"64",x"75",x"72",x"63",x"68",x"20",x"4E",x"75", -- 35D0-35DF 
  x"6C",x"6C",x"20",x"57",x"6F",x"72",x"74",x"20",x"6E",x"69",x"63",x"68",x"74",x"20",x"64",x"65", -- 35E0-35EF 
  x"66",x"69",x"6E",x"69",x"65",x"72",x"74",x"20",x"45",x"69",x"6E",x"67",x"61",x"62",x"65",x"7A", -- 35F0-35FF 
  x"65",x"69",x"6C",x"65",x"20",x"7A",x"75",x"20",x"6C",x"61",x"6E",x"67",x"20",x"53",x"74",x"72", -- 3600-360F 
  x"75",x"6B",x"74",x"75",x"72",x"66",x"65",x"68",x"6C",x"65",x"72",x"20",x"69",x"6E",x"20",x"49", -- 3610-361F 
  x"46",x"20",x"45",x"4E",x"44",x"5F",x"49",x"46",x"20",x"42",x"45",x"47",x"49",x"4E",x"20",x"55", -- 3620-362F 
  x"4E",x"54",x"49",x"4C",x"20",x"44",x"4F",x"20",x"4C",x"4F",x"4F",x"50",x"20",x"20",x"6E",x"65", -- 3630-363F 
  x"67",x"61",x"74",x"69",x"76",x"65",x"72",x"20",x"45",x"78",x"70",x"6F",x"6E",x"65",x"6E",x"74", -- 3640-364F 
  x"20",x"5A",x"61",x"68",x"6C",x"65",x"6E",x"73",x"70",x"65",x"69",x"63",x"68",x"65",x"72",x"20", -- 3650-365F 
  x"76",x"6F",x"6C",x"6C",x"20",x"67",x"72",x"6F",x"C3",x"9F",x"65",x"20",x"67",x"61",x"6E",x"7A", -- 3660-366F 
  x"65",x"20",x"5A",x"61",x"68",x"6C",x"65",x"6E",x"20",x"6B",x"6F",x"6D",x"70",x"69",x"6C",x"69", -- 3670-367F 
  x"65",x"72",x"65",x"6E",x"20",x"67",x"65",x"68",x"74",x"20",x"6D",x"6F",x"6D",x"65",x"6E",x"74", -- 3680-368F 
  x"61",x"6E",x"20",x"6E",x"69",x"63",x"68",x"74",x"2C",x"20",x"73",x"69",x"65",x"68",x"65",x"20", -- 3690-369F 
  x"54",x"45",x"53",x"54",x"46",x"55",x"45",x"52",x"4E",x"45",x"55",x"45",x"53",x"2E",x"54",x"58", -- 36A0-36AF 
  x"54",x"20",x"53",x"54",x"52",x"47",x"3A",x"20",x"5E",x"47",x"20",x"2F",x"31",x"78",x"50",x"49", -- 36B0-36BF 
  x"45",x"50",x"2F",x"20",x"5E",x"46",x"20",x"51",x"55",x"49",x"54",x"20",x"5E",x"41",x"20",x"41", -- 36C0-36CF 
  x"6E",x"67",x"65",x"68",x"61",x"6C",x"74",x"65",x"6E",x"20",x"66",x"C3",x"BC",x"72",x"20",x"67", -- 36D0-36DF 
  x"65",x"6E",x"61",x"75",x"20",x"65",x"69",x"6E",x"65",x"20",x"45",x"69",x"6E",x"67",x"61",x"62", -- 36E0-36EF 
  x"65",x"7A",x"65",x"69",x"6C",x"65",x"3A",x"20",x"20",x"6F",x"6B",x"20",x"51",x"55",x"45",x"52", -- 36F0-36FF 
  x"59",x"20",x"28",x"2A",x"52",x"45",x"4D",x"2A",x"29",x"20",x"2F",x"6F",x"6B",x"3E",x"20",x"28", -- 3700-370F 
  x"2A",x"45",x"4E",x"44",x"2A",x"29",x"20",x"6F",x"6B",x"3E",x"20",x"48",x"45",x"58",x"20",x"44", -- 3710-371F 
  x"45",x"43",x"49",x"4D",x"41",x"4C",x"20",x"4E",x"4C",x"49",x"54",x"2C",x"20",x"4D",x"2E",x"20", -- 3720-372F 
  x"4D",x"2B",x"20",x"4D",x"2D",x"20",x"4D",x"2A",x"20",x"4D",x"2F",x"20",x"4D",x"2F",x"4D",x"4F", -- 3730-373F 
  x"44",x"20",x"4D",x"4D",x"4F",x"44",x"20",x"2E",x"20",x"2B",x"20",x"2D",x"20",x"2A",x"20",x"2F", -- 3740-374F 
  x"20",x"2F",x"4D",x"4F",x"44",x"20",x"47",x"47",x"54",x"20",x"42",x"4B",x"20",x"5E",x"20",x"3F", -- 3750-375F 
  x"20",x"29",x"20",x"28",x"3A",x"29",x"20",x"49",x"4D",x"4D",x"45",x"44",x"49",x"41",x"54",x"45", -- 3760-376F 
  others=>x"00");

-- Rückkehrstapel
type stapRAMTYPE is array(0 to 1024-1) of STD_LOGIC_VECTOR (15 downto 0);
shared variable stapR: stapRAMTYPE:=(
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C00-2C0F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C10-2C1F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C20-2C2F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C30-2C3F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C40-2C4F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C50-2C5F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C60-2C6F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C70-2C7F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C80-2C8F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C90-2C9F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2CA0-2CAF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2CB0-2CBF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2CC0-2CCF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2CD0-2CDF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2CE0-2CEF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2CF0-2CFF 
  x"0000",x"0000",x"0000",x"0000",x"0055",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D00-2D0F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D10-2D1F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D20-2D2F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D30-2D3F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D40-2D4F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D50-2D5F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D60-2D6F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D70-2D7F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D80-2D8F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D90-2D9F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2DA0-2DAF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2DB0-2DBF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2DC0-2DCF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2DD0-2DDF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2DE0-2DEF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2DF0-2DFF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E00-2E0F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E10-2E1F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E20-2E2F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E30-2E3F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E40-2E4F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E50-2E5F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E60-2E6F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E70-2E7F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E80-2E8F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E90-2E9F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2EA0-2EAF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2EB0-2EBF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2EC0-2ECF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2ED0-2EDF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0008", -- 2EE0-2EEF 
  x"0008",x"0000",x"0001",x"2F1A",x"0000",x"0001",x"2F1B",x"1410",x"0008",x"3B0A",x"0001",x"0001",x"3B45",x"00BB",x"0001",x"FFFF", -- 2EF0-2EFF 
  x"0000",x"0000",x"3000",x"3F42",x"3F42",x"FFFF",x"3761",x"125E",x"0010",x"3B00",x"3B00",x"3B0C",x"3B12",x"3B45",x"0000",x"125E", -- 2F00-2F0F 
  x"0000",x"1257",x"3000",x"3761",x"0028",x"0062",x"0000",x"2F00",x"2F22",x"0000",x"0000",x"140C",x"1400",x"2000",x"0001",x"1400", -- 2F10-2F1F 
  x"1400",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F20-2F2F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F30-2F3F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F40-2F4F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F50-2F5F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F60-2F6F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F70-2F7F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F80-2F8F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F90-2F9F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2FA0-2FAF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2FB0-2FBF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2FC0-2FCF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0301",x"0301",x"0301",x"0301",x"0301",x"0301",x"0301",x"0301", -- 2FD0-2FDF 
  x"0301",x"0301",x"0301",x"0301",x"0446",x"02DB",x"0053",x"02A3",x"02DB",x"02DB",x"02DB",x"02DB",x"02DB",x"065F",x"02DB",x"0053", -- 2FE0-2FEF 
  x"02DB",x"02DB",x"02DB",x"0053",x"0322",x"0349",x"01FA",x"0296",x"081C",x"FFFF",x"06FB",x"3B05",x"3B06",x"3B00",x"3B00",x"0745", -- 2FF0-2FFF 
  others=>x"0000");

--diese Funktion übernimmt von SP nur die beiden niedrigsten Bits
  function P(SP : integer) return integer is begin
--    return CONV_INTEGER(CONV_UNSIGNED(SP,2));
    return SP mod 4;
    end;

-- alles Signale um die Stapel-RAM's zu machen.
signal HOLE_VOM_STAPEL,STORE_ZUM_STAPEL,ADRESSE_ZUM_STAPEL: REG;
signal WE_ZUM_STAPEL: STD_LOGIC_VECTOR (3 downto 0);
type STAPELTYPE is array(0 to 31) of STD_LOGIC_VECTOR (15 downto 0);
signal stap1,stap2,stap3,stap0: STAPELTYPE:=(others=>x"0000");
-- Rueckkehrstapel
signal RPC,RPCC: STD_LOGIC_VECTOR (15 downto 0);
signal RP: STD_LOGIC_VECTOR (15 downto 0):=x"3000";
signal RW: STD_LOGIC;
-- kompletten Speicher anschliessen
signal PC_ZUM_ProgRAM,PD_VOM_ProgRAM: STD_LOGIC_VECTOR (15 downto 0);
signal STORE_ZUM_RAM,EXFET,ADRESSE_ZUM_RAM: STD_LOGIC_VECTOR (15 downto 0);
signal FETCH_VOM_ProgRAM,FETCH_VOM_ByteRAM,FETCH_VOM_stapR: STD_LOGIC_VECTOR (15 downto 0);
signal WE_ZUM_RAM,WE_ZUM_ProgRAM,WE_ZUM_ByteRAM,WE_ZUM_stapR: STD_LOGIC;
-- fuer EMIT-Ausgabe
signal EMIT_ABGESCHICKT_LOCAL,EMIT_ANGEKOMMEN_RUHEND,XOFF_INPUT_L: STD_LOGIC:='0';
signal KEY_ANGEKOMMEN_LOCAL,KEY_ABGESCHICKT_RUHEND,KEY_ABGESCHICKT_MERK: STD_LOGIC:='0';
signal KEY_BYTE_RUHEND: STD_LOGIC_VECTOR (7 downto 0);


begin

process begin wait until (CLK_I'event and CLK_I='1'); --ruhende Eingangsdaten für FortyForthprocessor
  EMIT_ANGEKOMMEN_RUHEND<=EMIT_ANGEKOMMEN;
  KEY_BYTE_RUHEND<=KEY_BYTE;
  KEY_ABGESCHICKT_RUHEND<=KEY_ABGESCHICKT;
  end process;
  

process -- FortyForthProcessor
variable PC,PD,ADR,DAT,DIST: STD_LOGIC_VECTOR (15 downto 0):=x"0000";
variable WE: STD_LOGIC;
variable SP: integer:=0;
variable R: REG:=(others=>x"0000");
-- Stapeleintraege benennen
variable A,B,C,D: STD_LOGIC_VECTOR (15 downto 0):=x"0000";
variable T: integer range 0 to 4;
variable W: STD_LOGIC_VECTOR (3 downto 0);
-- fuer Umstapeln 
variable STAK: STD_LOGIC_VECTOR (7 downto 0);
-- fuer Rechenoperationen mit Uebertrag
variable U: STD_LOGIC_VECTOR (31 downto 0);
-- fuer Division
variable UBIT: STD_LOGIC;
-- fuer Supermult
variable SUMME: STD_LOGIC_VECTOR (31 downto 0);

begin wait until (CLK_I'event and CLK_I='0'); PC_SIM<=PC;--Simulation
  -- ob ein KEY aingetroffen ist --
  if KEY_ABGESCHICKT_MERK/=KEY_ABGESCHICKT_RUHEND then 
    KEY_ABGESCHICKT_MERK<=KEY_ABGESCHICKT_RUHEND;
    PD:=x"4026";
    PC:=PC;
    else
      PD:=PD_VOM_ProgRAM;
      PC:=PC+1;
      end if;                                           -- Simulation --
  WE:='0';                                              PD_SIM<=PD;
  DIST:=PD(11)&PD(11)&PD(11)&PD(11)&PD(11 downto 0);    SP_SIM<=SP;
  -- oberste 4 Stapeleintraege entnehmen
  R:=HOLE_VOM_STAPEL;                                   -- Simulation --
  A:=R(P(SP-1));                                        A_SIM<=A;
  B:=R(P(SP-2));                                        B_SIM<=B;
  C:=R(P(SP-3));                                        C_SIM<=C;
  D:=R(P(SP-4));                                        D_SIM<=D;
  T:=0;
  -- Rueckkehrstapel
  RW<='0';
 
  if PD(15 downto 13)="010" then                 -- 4000-5FFF Unterprogrammaufruf
    RPC<=PC;PC:=PD and x"3FFF";RP<=RP-1;RW<='1';
    elsif PD(15 downto 12)=x"8" then PC:=PC+DIST;-- 8000-8FFF relativer Sprung
    elsif PD(15 downto 12)=x"9" then             -- 9000-9FFF bedingter relativer Sprung
      if A=x"0000" then PC:=PC+DIST; end if; SP:=SP-1;
    elsif PD=x"A003" then PC:=RPCC;RP<=RP+1;     -- ; Rückkehr aus Unterprogramm
    elsif PD=x"A00D" then -- 0= Vergleich ob gleich Null
      if A=x"0000" then A:=x"FFFF"; 
        else A:=x"0000"; end if;
      T:=1;
    elsif PD=x"A00F" then -- 0< Vergleich ob kleiner Null
      if A>=x"8000" then A:=x"FFFF";
        else A:=x"0000"; end if;
      T:=1;
    elsif PD=x"A000" then -- MINUS Vorzeichen wechseln
      A:=(not A)+1;
      T:=1;
    elsif PD=x"A00B" then -- NOT Bitweises Komplement
      A:=not A;
      T:=1;
    elsif PD=x"A008" then -- AND Bitweises Und
      A:=B and A; 
      T:=1;
      SP:=SP-1;
    elsif PD=x"A00E" then -- OR Bitweises Oder
      A:=B or A; 
      T:=1;
      SP:=SP-1;
    elsif PD=x"A007" then -- + Addition
      A:=B+A; 
      T:=1;
      SP:=SP-1;
    elsif PD=x"A001" then -- U+ Addition mit Übertrag
      U:=(x"0000"&C)+(x"0000"&B)+(x"0000"&A);
      B:=U(31 downto 16);
      A:=U(15 downto 0);
      T:=2;
      SP:=SP-1;
    elsif PD=x"A002" then -- U* Multiplikation mit Übertrag
      U:=(x"0000"&C)+B*A;
      B:=U(31 downto 16);
      A:=U(15 downto 0);
      T:=2;
      SP:=SP-1;
    elsif PD=x"A005" then -- EMIT Zeichen ausgeben
      if (EMIT_ABGESCHICKT_LOCAL=EMIT_ANGEKOMMEN_RUHEND) and XOFF_INPUT_L='0' then
        EMIT_BYTE<=A(7 downto 0);
        EMIT_ABGESCHICKT_LOCAL<=not EMIT_ANGEKOMMEN_RUHEND;
        T:=0;
        SP:=SP-1;
        else PC:=PC-1; end if; -- warten
    elsif PD=x"A009" then -- STORE Speicheradresse beschreiben
      case A is
        when x"2800" => KEY_ANGEKOMMEN_LOCAL<=not KEY_ANGEKOMMEN_LOCAL;
        when x"2801" => SP:=CONV_INTEGER(B);
        when x"2802" => RP<=B;
        when x"2803" => PC:=B;
        when others => ADR:=A;DAT:=B;WE:='1' ;
        end case;
      T:=0;
      SP:=SP-2;
    elsif PD=x"A00A" then -- FETCH Speicheradresse lesen
      case A is
        when x"2800" => A:=x"00"&KEY_BYTE_RUHEND;
        when x"2801" => A:=CONV_STD_LOGIC_VECTOR(SP-1,16);
        when x"2802" => A:=RP;
        when x"2803" => A:=PC;
        when others => A:=EXFET;
        end case;
      T:=1;
    elsif PD=x"A014" then -- DI32 DIVISION_MIT_REST 32B/16B=16R/16Q
      UBIT:=C(15);
      C:=C(14 downto 0)&B(15);
      B:=B(14 downto 0)&'0';
      if (UBIT&C)>=('0'&A) then
        C:=C-A;
        B(0):='1';
        end if;
      T:=3;
    elsif PD=x"A017" then -- MULT_I
      --     D    C    B    A        stapR
      --     c    ü   adr1 adr2      i
      -- c   ü   erg1 adr2 adr1      i-1
      SUMME:=(D*EXFET)+(x"0000"&C);
      C:=A;A:=B;B:=C;
      D:=SUMME(31 downto 16); 
      C:=SUMME(15 downto 0);
      RPC<=RPCC-1; RW<='1';
      T:=4; SP:=SP+1;
    elsif PD=x"A018" then -- MULT_II
      --     D    C     B      A         stapR
      -- c   ü1  erg1   adr2   adr1      i-1
      -- c   ü2  adr1+1 adr2+1 i-1       i-1
      SUMME:=(D&C)+(x"0000"&EXFET);
      D:=SUMME(31 downto 16); 
      DAT:=SUMME(15 downto 0);
      ADR:=A;
      WE:='1';
      C:=A+1;
      B:=B+1;
      if RPCC=x"0000" then A:=x"FFFF"; else A:=x"0000"; end if;
      T:=4;
    elsif PD(15 downto 12)=x"B" then           -- B000-BFFF Umstapeln
      STAK:="00000000";
      if PD(7)='1' then STAK:=STAK(5 downto 0)&"11"; T:=T+1; end if;
      if PD(6)='1' then STAK:=STAK(5 downto 0)&"10"; T:=T+1; end if;
      if PD(5)='1' then STAK:=STAK(5 downto 0)&"01"; T:=T+1; end if;
      if PD(4)='1' then STAK:=STAK(5 downto 0)&"00"; T:=T+1; end if;
      if PD(3)='1' then STAK:=STAK(5 downto 0)&"11"; T:=T+1; end if;
      if PD(2)='1' then STAK:=STAK(5 downto 0)&"10"; T:=T+1; end if;
      if PD(1)='1' then STAK:=STAK(5 downto 0)&"01"; T:=T+1; end if;
      if PD(0)='1' then STAK:=STAK(5 downto 0)&"00"; T:=T+1; end if;
      A:=R(P(SP-1-CONV_INTEGER(STAK(1 downto 0))));
      B:=R(P(SP-1-CONV_INTEGER(STAK(3 downto 2))));
      C:=R(P(SP-1-CONV_INTEGER(STAK(5 downto 4))));
      D:=R(P(SP-1-CONV_INTEGER(STAK(7 downto 6))));
      SP:=SP+CONV_INTEGER(PD(11 downto 8))-4;
    else A:=PD; SP:=SP+1; T:=1; end if;                    -- LIT
    
  -- oberste T Stapeleintraege zurückspeichern
  W:="0000";
  if T/=0 then R(P(SP-1)):=A; W(P(SP-1)):='1';
    if T/=1 then R(P(SP-2)):=B; W(P(SP-2)):='1';
      if T/=2 then R(P(SP-3)):=C; W(P(SP-3)):='1';
        if T/=3 then R(P(SP-4)):=D; W(P(SP-4)):='1';
          end if; end if; end if; end if;
  -- Ausgabeadresse zum StapRAM zusammenbasteln
  ADRESSE_ZUM_STAPEL(0)<=CONV_STD_LOGIC_VECTOR(SP-1,16);
  ADRESSE_ZUM_STAPEL(1)<=CONV_STD_LOGIC_VECTOR(SP-2,16);
  ADRESSE_ZUM_STAPEL(2)<=CONV_STD_LOGIC_VECTOR(SP-3,16);
  ADRESSE_ZUM_STAPEL(3)<=CONV_STD_LOGIC_VECTOR(SP-4,16);
  STORE_ZUM_STAPEL<=R;
  WE_ZUM_STAPEL<=W;
  -- ADR, DAT, WE, PC
  if WE='1' then ADRESSE_ZUM_RAM<=ADR; else ADRESSE_ZUM_RAM<=R(P(SP-1)); end if;
  STORE_ZUM_RAM<=DAT;
  WE_ZUM_RAM<=WE;
  PC_ZUM_ProgRAM<=PC;
  end process;

ADR_O<=ADRESSE_ZUM_RAM;
DAT_O<=STORE_ZUM_RAM;
WE_O<=WE_ZUM_RAM;
EMIT_ABGESCHICKT<=EMIT_ABGESCHICKT_LOCAL;
KEY_ANGEKOMMEN<=KEY_ANGEKOMMEN_LOCAL;

-- hier werden die Lesedaten der unterschiedlichen Speicher zusammengefuehrt
EXFET<=FETCH_VOM_ProgRAM when ADRESSE_ZUM_RAM(15 downto 13)="000" else
       FETCH_VOM_stapR when ADRESSE_ZUM_RAM(15 downto 10)="001011" else
       x"00"&FETCH_VOM_ByteRAM(7 downto 0) when ADRESSE_ZUM_RAM(15 downto 12)="0011" else
       DAT_I;

-- hier wird WE auf die unterschiedlichen Speicher aufgeteilt
WE_ZUM_ProgRAM<=WE_ZUM_RAM when ADRESSE_ZUM_RAM(15 downto 13)="000" else '0';
WE_ZUM_stapR  <=WE_ZUM_RAM when ADRESSE_ZUM_RAM(15 downto 10)="001011" else '0';
WE_ZUM_ByteRAM<=WE_ZUM_RAM when ADRESSE_ZUM_RAM(15 downto 12)="0011" else '0';


process -- Programmspeicher 0000H-1FFFH,
begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_ProgRAM='1' then 
    ProgRAM(CONV_INTEGER(ADRESSE_ZUM_RAM(12 downto 0)))<=STORE_ZUM_RAM; 
    FETCH_VOM_ProgRAM<=STORE_ZUM_RAM; 
	  else
      FETCH_VOM_ProgRAM<=ProgRAM(CONV_INTEGER(ADRESSE_ZUM_RAM(12 downto 0)));
      end if;
  PD_VOM_ProgRAM<=ProgRAM(CONV_INTEGER(PC_ZUM_ProgRAM(12 downto 0)));
  end process;

process -- Textspeicher 3000H-3FFFH
begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_ByteRAM='1' then 
    ByteRAM(CONV_INTEGER(ADRESSE_ZUM_RAM(12 downto 0)))<=STORE_ZUM_RAM(7 downto 0); 
    FETCH_VOM_ByteRAM<=STORE_ZUM_RAM; 
	 else
      FETCH_VOM_ByteRAM<=x"00"&ByteRAM(CONV_INTEGER(ADRESSE_ZUM_RAM(12 downto 0)));
      end if;
  end process;

process --Rueckkehrstapel, TRUE_DUAL_PORT
begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_StapR='1' then 
    stapR(CONV_INTEGER(ADRESSE_ZUM_RAM(9 downto 0))):=STORE_ZUM_RAM; 
    end if;
  FETCH_VOM_stapR<=stapR(CONV_INTEGER(ADRESSE_ZUM_RAM(9 downto 0)));
  end process;
process begin wait until (CLK_I'event and CLK_I='1');
  if RW='1' then
    stapR(CONV_INTEGER(RP(9 downto 0))):=RPC;
    RPCC<=RPC;
     else
      RPCC<=stapR(CONV_INTEGER(RP(9 downto 0)));
    end if;
  end process;

--StapelRAM:
process begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_STAPEL(0)='1' then
    stap0(CONV_INTEGER(ADRESSE_ZUM_STAPEL(0)(6 downto 2)))<=STORE_ZUM_STAPEL(0);
    HOLE_VOM_STAPEL(0)<=STORE_ZUM_STAPEL(0);
     else
      HOLE_VOM_STAPEL(0)<=stap0(CONV_INTEGER(ADRESSE_ZUM_STAPEL(0)(6 downto 2)));
    end if;
  end process;
process begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_STAPEL(1)='1' then
    stap1(CONV_INTEGER(ADRESSE_ZUM_STAPEL(1)(6 downto 2)))<=STORE_ZUM_STAPEL(1);
    HOLE_VOM_STAPEL(1)<=STORE_ZUM_STAPEL(1);
     else
      HOLE_VOM_STAPEL(1)<=stap1(CONV_INTEGER(ADRESSE_ZUM_STAPEL(1)(6 downto 2)));
    end if;
  end process;
process begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_STAPEL(2)='1' then
    stap2(CONV_INTEGER(ADRESSE_ZUM_STAPEL(2)(6 downto 2)))<=STORE_ZUM_STAPEL(2);
    HOLE_VOM_STAPEL(2)<=STORE_ZUM_STAPEL(2);
     else
      HOLE_VOM_STAPEL(2)<=stap2(CONV_INTEGER(ADRESSE_ZUM_STAPEL(2)(6 downto 2)));
    end if;
  end process;
process begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_STAPEL(3)='1' then
    stap3(CONV_INTEGER(ADRESSE_ZUM_STAPEL(3)(6 downto 2)))<=STORE_ZUM_STAPEL(3);
    HOLE_VOM_STAPEL(3)<=STORE_ZUM_STAPEL(3);
     else
      HOLE_VOM_STAPEL(3)<=stap3(CONV_INTEGER(ADRESSE_ZUM_STAPEL(3)(6 downto 2)));
    end if;
  end process;

end Step_9;
