library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity FortyForthProcessor is
  Port (
    CLK_I: in STD_LOGIC;
    DAT_I: in STD_LOGIC_VECTOR (15 downto 0);
    ADR_O: out STD_LOGIC_VECTOR (15 downto 0);
    DAT_O: out STD_LOGIC_VECTOR (15 downto 0);
    WE_O: out STD_LOGIC;
    
    -- EMIT --
    EMIT_ABGESCHICKT: out STD_LOGIC;
    EMIT_BYTE: out STD_LOGIC_VECTOR (7 downto 0);
    EMIT_ANGEKOMMEN: in STD_LOGIC;
    
     -- EMIT --
    KEY_ABGESCHICKT: in STD_LOGIC;
    KEY_BYTE: in STD_LOGIC_VECTOR (7 downto 0);
    KEY_ANGEKOMMEN: out STD_LOGIC;

   -- nur zur Simulation und Fehlersuche:
    PC_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    PD_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    SP_SIM: out integer;
    A_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    B_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    C_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    D_SIM: out STD_LOGIC_VECTOR (15 downto 0)
    );
end FortyForthProcessor;

architecture Step_9 of FortyForthProcessor is

type REG is array(0 to 3) of STD_LOGIC_VECTOR (15 downto 0);
type RAMTYPE is array(0 to 8*1024-1) of STD_LOGIC_VECTOR (15 downto 0);
-- Programmspeicher 0000H-1FFFH
signal ProgRAM: RAMTYPE:=(
  x"4010",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 0000-000F 
  x"479C",x"A003",x"44E9",x"9001",x"A003",x"B300",x"8000",x"8FFA",x"0000",x"111C",x"0000",x"0000",x"0000",x"0000",x"1111",x"1107", -- 0010-001F 
  x"4000",x"A003",x"4000",x"A003",x"4000",x"A003",x"44BA",x"A003",x"4000",x"A003",x"4000",x"A003",x"4000",x"A003",x"4000",x"A003", -- 0020-002F 
  x"4000",x"A003",x"4000",x"A003",x"4000",x"A003",x"4000",x"A003",x"4000",x"A003",x"4000",x"A003",x"4000",x"A003",x"4000",x"A003", -- 0030-003F 
--                --RP0--
  x"0000",x"0000",x"4000",x"FC73",x"FC73",x"FFFF",x"E72D",x"11D6",x"0010",x"FB00",x"FB00",x"FB09",x"FB0F",x"FB45",x"0000",x"11D6", -- 0040-004F 
  x"0000",x"11CF",x"E000",x"E72D",x"0058",x"0049",x"0000",x"2FEF",x"0000",x"E000",x"0001",x"47AF",x"0029",x"4621",x"B200",x"A003", -- 0050-005F 
  x"FFF8",x"E002",x"0001",x"47AF",x"0000",x"0050",x"A009",x"A003",x"FFF8",x"E004",x"0001",x"47BD",x"0001",x"0050",x"A009",x"A003", -- 0060-006F 
  x"FFF8",x"E006",x"0007",x"47AF",x"0020",x"4621",x"469B",x"46DB",x"B300",x"46E4",x"A003",x"FFF5",x"E00E",x"0006",x"47B6",x"42FA", -- 0070-007F 
  x"B501",x"42AD",x"430D",x"A00A",x"A003",x"FFF6",x"E015",x"0004",x"47BD",x"5167",x"A003",x"42D4",x"B502",x"C000",x"42C2",x"A00E", -- 0080-008F 
  x"9001",x"407E",x"432D",x"A003",x"FFF1",x"E01A",x"000B",x"47B6",x"42FA",x"A00A",x"0050",x"A00A",x"9001",x"4089",x"A003",x"FFF5", -- 0090-009F 
  x"E026",x"0008",x"47BD",x"46ED",x"4097",x"432D",x"47A7",x"A003",x"FFF7",x"E02F",x"0002",x"4098",x"D001",x"FFFB",x"E032",x"0002", -- 00A0-00AF 
  x"4098",x"D002",x"FFFB",x"E035",x"0002",x"4098",x"D003",x"FFFB",x"E038",x"0004",x"4098",x"0040",x"FFFB",x"E03D",x"0009",x"4098", -- 00B0-00BF 
  x"0041",x"FFFB",x"E047",x"0003",x"4098",x"0042",x"FFFB",x"E04B",x"0007",x"4098",x"0043",x"FFFB",x"E053",x"0007",x"4098",x"0044", -- 00C0-00CF 
  x"FFFB",x"E05B",x"0004",x"4098",x"0045",x"FFFB",x"E060",x"0007",x"4098",x"0046",x"FFFB",x"E068",x"0004",x"4098",x"0047",x"FFFB", -- 00D0-00DF 
  x"E06D",x"0004",x"4098",x"0048",x"FFFB",x"E072",x"0003",x"4098",x"0049",x"FFFB",x"E076",x"0003",x"4098",x"004A",x"FFFB",x"E07A", -- 00E0-00EF 
  x"0003",x"4098",x"004B",x"FFFB",x"E07E",x"0003",x"4098",x"004C",x"FFFB",x"E082",x"0003",x"4098",x"004D",x"FFFB",x"E086",x"0007", -- 00F0-00FF 
  x"4098",x"004E",x"FFFB",x"E08E",x"0002",x"4098",x"004F",x"FFFB",x"E091",x"0004",x"4098",x"0050",x"FFFB",x"E096",x"0003",x"4098", -- 0100-010F 
  x"0051",x"FFFB",x"E09A",x"0004",x"4098",x"0052",x"FFFB",x"E09F",x"0005",x"4098",x"0053",x"FFFB",x"E0A5",x"0006",x"4098",x"0054", -- 0110-011F 
  x"FFFB",x"E0AC",x"0003",x"4098",x"0055",x"FFFB",x"E0B0",x"0009",x"4098",x"0056",x"FFFB",x"E0BA",x"0007",x"4098",x"01AC",x"FFFB", -- 0120-012F 
  x"E0C2",x"0006",x"4098",x"A003",x"FFFB",x"E0C9",x"0008",x"47B6",x"42FA",x"0050",x"A00A",x"9003",x"A00A",x"432D",x"8001",x"4338", -- 0130-013F 
  x"A003",x"FFF3",x"E0D2",x"0005",x"47BD",x"46ED",x"4137",x"432D",x"407F",x"A003",x"432D",x"47A7",x"A003",x"FFF4",x"E0D8",x"0005", -- 0140-014F 
  x"4138",x"A000",x"A003",x"FFFA",x"E0DE",x"0002",x"4138",x"A001",x"A003",x"FFFA",x"E0E1",x"0002",x"4138",x"A002",x"A003",x"FFFA", -- 0150-015F 
  x"E0E4",x"0002",x"4138",x"A00D",x"A003",x"FFFA",x"E0E7",x"0003",x"4138",x"A00F",x"A003",x"FFFA",x"E0EB",x"0008",x"4138",x"A005", -- 0160-016F 
  x"A003",x"FFFA",x"E0F4",x"0003",x"4138",x"A00B",x"A003",x"FFFA",x"E0F8",x"0003",x"4138",x"A008",x"A003",x"FFFA",x"E0FC",x"0002", -- 0170-017F 
  x"4138",x"A00E",x"A003",x"FFFA",x"E0FF",x"0007",x"4138",x"A00C",x"A003",x"FFFA",x"E107",x"0001",x"4138",x"A007",x"A003",x"FFFA", -- 0180-018F 
  x"E109",x"0001",x"4138",x"A009",x"A003",x"FFFA",x"E10B",x"0001",x"4138",x"A00A",x"A003",x"FFFA",x"E10D",x"0004",x"4138",x"B412", -- 0190-019F 
  x"A003",x"FFFA",x"E112",x"0004",x"4138",x"B502",x"A003",x"FFFA",x"E117",x"0003",x"4138",x"B501",x"A003",x"FFFA",x"E11B",x"0003", -- 01A0-01AF 
  x"4138",x"B434",x"A003",x"FFFA",x"E11F",x"0004",x"4138",x"B300",x"A003",x"FFFA",x"E124",x"0005",x"4138",x"B43C",x"A003",x"FFFA", -- 01B0-01BF 
  x"E12A",x"0005",x"4138",x"B60C",x"A003",x"FFFA",x"E130",x"0004",x"4138",x"B603",x"A003",x"FFFA",x"E135",x"0005",x"4138",x"B200", -- 01C0-01CF 
  x"A003",x"FFFA",x"E13B",x"0004",x"4138",x"8000",x"A003",x"FFFA",x"E140",x"0002",x"47BD",x"0053",x"A00A",x"A009",x"0001",x"0053", -- 01D0-01DF 
  x"42EF",x"A003",x"FFF5",x"E143",x"0002",x"47BD",x"0053",x"A00A",x"4089",x"B501",x"432D",x"B412",x"B501",x"A00A",x"41DB",x"42AD", -- 01E0-01EF 
  x"B412",x"0001",x"42B4",x"B501",x"A00D",x"9FF5",x"B200",x"0020",x"41DB",x"A003",x"FFE8",x"E146",x"0007",x"47B6",x"4621",x"0050", -- 01F0-01FF 
  x"A00A",x"9003",x"41E6",x"42FA",x"46E4",x"A003",x"FFF4",x"E14E",x"0005",x"47BD",x"46ED",x"0001",x"0050",x"A009",x"432D",x"41FD", -- 0200-020F 
  x"FFFF",x"0055",x"42EF",x"A003",x"FFF2",x"E154",x"0001",x"0022",x"41FE",x"A003",x"FFFA",x"E156",x"0002",x"0022",x"41FE",x"4365", -- 0210-021F 
  x"A003",x"FFF9",x"E159",x"0004",x"47BD",x"004F",x"A00A",x"A003",x"FFF9",x"E15E",x"0005",x"47BD",x"0008",x"A003",x"FFFA",x"E164", -- 0220-022F 
  x"0006",x"47BD",x"0009",x"A003",x"FFFA",x"E16B",x"0006",x"47BD",x"1000",x"42DB",x"B412",x"0FFF",x"A008",x"A00E",x"A003",x"FFF5", -- 0230-023F 
  x"E172",x"0005",x"47BD",x"004F",x"42EF",x"A003",x"FFF9",x"E178",x"0007",x"47BD",x"4225",x"42AD",x"42B4",x"422C",x"4238",x"432D", -- 0240-024F 
  x"A003",x"FFF5",x"E180",x"0008",x"47BD",x"4225",x"42AD",x"42B4",x"4232",x"4238",x"432D",x"A003",x"FFF5",x"E189",x"0005",x"47AF", -- 0250-025F 
  x"4225",x"A003",x"FFFA",x"E18F",x"0005",x"47AF",x"424A",x"A003",x"FFFA",x"E195",x"0005",x"47AF",x"4255",x"A003",x"FFFA",x"E19B", -- 0260-026F 
  x"0002",x"47AF",x"4232",x"0001",x"4243",x"4225",x"A003",x"FFF7",x"E19E",x"0006",x"47AF",x"4225",x"B502",x"42B4",x"B434",x"4238", -- 0270-027F 
  x"B412",x"0001",x"42B4",x"A009",x"A003",x"FFF2",x"E1A5",x"0004",x"47AF",x"0001",x"4243",x"427A",x"422C",x"4225",x"A003",x"FFF6", -- 0280-028F 
  x"E1AA",x"0005",x"47AF",x"4271",x"A003",x"FFFA",x"E1B0",x"0006",x"47AF",x"B434",x"4265",x"427A",x"A003",x"FFF8",x"E1B7",x"0002", -- 0290-029F 
  x"47BD",x"A00A",x"A003",x"FFFA",x"E1BA",x"0002",x"47BD",x"A009",x"A003",x"FFFA",x"E1BD",x"0002",x"47BD",x"0001",x"A007",x"A003", -- 02A0-02AF 
  x"FFF9",x"E1C0",x"0001",x"47BD",x"A000",x"A007",x"A003",x"FFF9",x"E1C2",x"0001",x"47BD",x"42B4",x"A00D",x"A003",x"FFF9",x"E1C4", -- 02B0-02BF 
  x"0002",x"47BD",x"407F",x"8000",x"A007",x"B412",x"A00B",x"407F",x"8000",x"A007",x"0000",x"A001",x"B300",x"A00D",x"A00B",x"A003", -- 02C0-02CF 
  x"FFEE",x"E1C7",x"0001",x"47BD",x"B412",x"42C2",x"A003",x"FFF9",x"E1C9",x"0001",x"47BD",x"0000",x"B434",x"B434",x"A002",x"B412", -- 02D0-02DF 
  x"B300",x"A003",x"FFF5",x"E1CB",x"0003",x"47BD",x"E1CF",x"0004",x"421F",x"8FFC",x"A003",x"FFF7",x"E1D4",x"0002",x"47BD",x"B412", -- 02E0-02EF 
  x"B502",x"A00A",x"A007",x"B412",x"A009",x"A003",x"FFF5",x"E1D7",x"0002",x"47BD",x"D002",x"A00A",x"42AD",x"A00A",x"D002",x"A00A", -- 02F0-02FF 
  x"42AD",x"D002",x"B603",x"A00A",x"A00A",x"B412",x"A009",x"A009",x"A003",x"FFED",x"E1DA",x"0002",x"47BD",x"D002",x"A00A",x"B501", -- 0300-030F 
  x"FFFF",x"A007",x"D002",x"B603",x"A00A",x"A00A",x"B412",x"B501",x"FFFF",x"A007",x"D002",x"A009",x"A009",x"A009",x"A009",x"A003", -- 0310-031F 
  x"FFE9",x"E1DD",x"0001",x"47BD",x"D002",x"A00A",x"42AD",x"A00A",x"A003",x"FFF7",x"E1DF",x"0001",x"47BD",x"004F",x"A00A",x"A009", -- 0320-032F 
  x"0001",x"004F",x"42EF",x"A003",x"FFF5",x"E1E1",x"0007",x"47BD",x"D003",x"A009",x"A003",x"FFF9",x"E1E9",x"0003",x"47BD",x"0012", -- 0330-033F 
  x"4338",x"A003",x"FFF9",x"E1ED",x"0004",x"47BD",x"016F",x"4338",x"A003",x"FFF9",x"E1F2",x"0005",x"47BD",x"0000",x"B412",x"0010", -- 0340-034F 
  x"A002",x"B412",x"A003",x"FFF6",x"E1F8",x"0003",x"47BD",x"B501",x"000A",x"42C2",x"9001",x"8002",x"0007",x"A007",x"0030",x"A007", -- 0350-035F 
  x"A003",x"FFF2",x"E1FC",x"0004",x"47BD",x"B501",x"9009",x"B412",x"B501",x"42A1",x"4346",x"42AD",x"B412",x"0001",x"42B4",x"8FF5", -- 0360-036F 
  x"B200",x"A003",x"FFEF",x"E201",x"0003",x"47BD",x"434D",x"4357",x"4346",x"434D",x"4357",x"4346",x"434D",x"4357",x"4346",x"434D", -- 0370-037F 
  x"4357",x"4346",x"B300",x"A003",x"FFEE",x"E205",x"0002",x"47BD",x"4376",x"0020",x"4346",x"A003",x"FFF8",x"E208",x"0001",x"47BD", -- 0380-038F 
  x"4388",x"A003",x"FFFA",x"E20A",x"0001",x"47BD",x"A00A",x"4390",x"A003",x"FFF9",x"E20C",x"0002",x"47BD",x"0047",x"A00A",x"004F", -- 0390-039F 
  x"A00A",x"42B4",x"0050",x"A00A",x"A00D",x"A00B",x"A00E",x"0040",x"A00A",x"A00D",x"A00B",x"A008",x"9028",x"003C",x"4346",x"E20F", -- 03A0-03AF 
  x"0003",x"421F",x"0047",x"A00A",x"4390",x"0046",x"A00A",x"4390",x"003C",x"4346",x"E213",x"0004",x"421F",x"003C",x"4346",x"E218", -- 03B0-03BF 
  x"0003",x"421F",x"004F",x"A00A",x"4390",x"0053",x"A00A",x"4390",x"003C",x"4346",x"E21C",x"0004",x"421F",x"004F",x"A00A",x"0047", -- 03C0-03CF 
  x"A009",x"0053",x"A00A",x"0046",x"A009",x"000A",x"4346",x"A003",x"FFC1",x"E221",x"000A",x"47BD",x"A003",x"FFFB",x"E22C",x"0007", -- 03D0-03DF 
  x"47BD",x"439D",x"E234",x"0019",x"421F",x"0020",x"4346",x"0008",x"4346",x"433F",x"001B",x"42BB",x"9FF8",x"A003",x"FFEF",x"E24E", -- 03E0-03EF 
  x"0005",x"47BD",x"B501",x"004E",x"A009",x"0000",x"0050",x"A009",x"439D",x"004A",x"A00A",x"004C",x"A00A",x"004A",x"A00A",x"42B4", -- 03F0-03FF 
  x"0001",x"42B4",x"4365",x"E254",x"0003",x"421F",x"E258",x"000A",x"4219",x"4702",x"439D",x"E263",x"0016",x"421F",x"4390",x"43E1", -- 0400-040F 
  x"474F",x"A003",x"FFDC",x"E27A",x"0004",x"47BD",x"D001",x"A00A",x"0055",x"A009",x"A003",x"FFF7",x"E27F",x"0004",x"47BD",x"D001", -- 0410-041F 
  x"A00A",x"0055",x"A00A",x"42B4",x"9002",x"0009",x"43F2",x"A003",x"FFF3",x"E284",x"0005",x"47BD",x"42FA",x"B412",x"B501",x"A000", -- 0420-042F 
  x"D002",x"A00A",x"A007",x"D002",x"A009",x"D002",x"A00A",x"0056",x"A00A",x"430D",x"0056",x"A009",x"430D",x"430D",x"A003",x"FFE9", -- 0430-043F 
  x"E28A",x"0009",x"47BD",x"42FA",x"42FA",x"42FA",x"0056",x"A009",x"D002",x"A00A",x"A007",x"D002",x"A009",x"430D",x"A003",x"FFF0", -- 0440-044F 
  x"E294",x"0002",x"47BD",x"0056",x"A00A",x"A003",x"FFF9",x"E297",x"0002",x"47BD",x"0056",x"A00A",x"42AD",x"A003",x"FFF8",x"E29A", -- 0450-045F 
  x"0002",x"47BD",x"0056",x"A00A",x"0002",x"A007",x"A003",x"FFF7",x"E29D",x"0002",x"47BD",x"0056",x"A00A",x"0003",x"A007",x"A003", -- 0460-046F 
  x"FFF7",x"E2A0",x"0002",x"47BD",x"0056",x"A00A",x"0004",x"A007",x"A003",x"FFF7",x"E2A3",x"0002",x"47BD",x"0056",x"A00A",x"0005", -- 0470-047F 
  x"A007",x"A003",x"FFF7",x"E2A6",x"0002",x"47BD",x"0056",x"A00A",x"0006",x"A007",x"A003",x"FFF7",x"E2A9",x"0002",x"47BD",x"0056", -- 0480-048F 
  x"A00A",x"0007",x"A007",x"A003",x"FFF7",x"E2AC",x"0001",x"47AF",x"0020",x"4621",x"469B",x"46DB",x"B300",x"42AD",x"0050",x"A00A", -- 0490-049F 
  x"9001",x"4089",x"A003",x"FFF1",x"E2AE",x"0005",x"47BD",x"B501",x"A00A",x"0001",x"A007",x"B501",x"03FF",x"A008",x"0000",x"42BB", -- 04A0-04AF 
  x"9002",x"0400",x"42B4",x"B412",x"A009",x"A003",x"FFED",x"E2B4",x"0007",x"47BD",x"D000",x"A00A",x"B501",x"0008",x"42C2",x"9009", -- 04B0-04BF 
  x"0018",x"A007",x"A00A",x"B501",x"9002",x"B501",x"4338",x"B300",x"8018",x"0043",x"A00A",x"A009",x"0043",x"44A7",x"0043",x"A00A", -- 04C0-04CF 
  x"0044",x"A00A",x"42B4",x"03FF",x"A008",x"0100",x"42D4",x"9009",x"0045",x"A00A",x"A00D",x"9005",x"FFFF",x"0045",x"A009",x"0013", -- 04D0-04DF 
  x"4346",x"0000",x"D000",x"A009",x"A003",x"FFD1",x"E2BC",x"0008",x"47BD",x"0044",x"A00A",x"0043",x"A00A",x"42BB",x"9003",x"0000", -- 04E0-04EF 
  x"0000",x"8018",x"0044",x"A00A",x"A00A",x"FFFF",x"0044",x"44A7",x"0043",x"A00A",x"0044",x"A00A",x"42B4",x"03FF",x"A008",x"0080", -- 04F0-04FF 
  x"42C2",x"9008",x"0045",x"A00A",x"9005",x"0000",x"0045",x"A009",x"0011",x"4346",x"A003",x"FFDA",x"E2C5",x"0006",x"47BD",x"0005", -- 0500-050F 
  x"442C",x"4462",x"A009",x"445A",x"A009",x"445A",x"A00A",x"4474",x"A009",x"433F",x"B501",x"0014",x"42BB",x"9004",x"B300",x"445A", -- 0510-051F 
  x"A00A",x"42A1",x"B501",x"007F",x"42BB",x"9002",x"B300",x"0008",x"B501",x"0008",x"42BB",x"9012",x"4474",x"A00A",x"445A",x"A00A", -- 0520-052F 
  x"42C2",x"900C",x"FFFF",x"445A",x"42EF",x"0001",x"4462",x"42EF",x"0008",x"4346",x"0020",x"4346",x"0008",x"4346",x"B501",x"0020", -- 0530-053F 
  x"42C2",x"9001",x"8012",x"FFFF",x"4462",x"42EF",x"4462",x"A00A",x"A00F",x"9002",x"0006",x"43F2",x"B501",x"4346",x"B501",x"445A", -- 0540-054F 
  x"A00A",x"42A7",x"0001",x"445A",x"42EF",x"B501",x"0020",x"42C2",x"B502",x"0008",x"42BB",x"A00B",x"A008",x"B412",x"001B",x"42BB", -- 0550-055F 
  x"A00B",x"A008",x"4462",x"A00A",x"A00D",x"A00E",x"9FB2",x"0020",x"4346",x"4474",x"A00A",x"445A",x"A00A",x"4474",x"A00A",x"42B4", -- 0560-056F 
  x"B603",x"A007",x"0000",x"B412",x"42A7",x"4443",x"A003",x"FF94",x"E2CC",x"0005",x"47BD",x"B501",x"0030",x"42C2",x"A00B",x"B502", -- 0570-057F 
  x"003A",x"42C2",x"A008",x"B502",x"0041",x"42C2",x"A00B",x"A00E",x"B501",x"9015",x"B412",x"0030",x"42B4",x"B501",x"000A",x"42C2", -- 0580-058F 
  x"A00B",x"9002",x"0007",x"42B4",x"B501",x"0048",x"A00A",x"42C2",x"A00B",x"9004",x"B300",x"B300",x"0000",x"0000",x"B412",x"A003", -- 0590-059F 
  x"FFD7",x"E2D2",x"0006",x"47BD",x"5169",x"A003",x"445A",x"A009",x"4453",x"A009",x"0000",x"445A",x"A00A",x"9063",x"B501",x"4462", -- 05A0-05AF 
  x"A009",x"0001",x"447D",x"A009",x"FFFF",x"4486",x"A009",x"4453",x"A00A",x"4462",x"A00A",x"A007",x"42A1",x"002B",x"42BB",x"9009", -- 05B0-05BF 
  x"4462",x"A00A",x"42AD",x"4462",x"A009",x"0000",x"4486",x"A009",x"8016",x"4453",x"A00A",x"4462",x"A00A",x"A007",x"42A1",x"002D", -- 05C0-05CF 
  x"42BB",x"900D",x"4462",x"A00A",x"42AD",x"4462",x"A009",x"0000",x"4486",x"A009",x"447D",x"A00A",x"A000",x"447D",x"A009",x"4486", -- 05D0-05DF 
  x"A00A",x"9FD2",x"4462",x"A00A",x"445A",x"A00A",x"42C2",x"9029",x"4453",x"A00A",x"4462",x"A00A",x"A007",x"42A1",x"B501",x"9015", -- 05E0-05EF 
  x"457B",x"A00B",x"9007",x"B300",x"445A",x"A00A",x"A000",x"445A",x"A009",x"800A",x"B412",x"0048",x"A00A",x"42DB",x"A007",x"4462", -- 05F0-05FF 
  x"A00A",x"42AD",x"4462",x"A009",x"8005",x"B300",x"4462",x"A00A",x"445A",x"A009",x"4462",x"A00A",x"445A",x"A00A",x"42C2",x"A00B", -- 0600-060F 
  x"9FD7",x"447D",x"A00A",x"A00F",x"9001",x"A000",x"4462",x"A00A",x"445A",x"A00A",x"42B4",x"4443",x"A003",x"FF83",x"E2D9",x"0004", -- 0610-061F 
  x"47BD",x"430D",x"004C",x"A00A",x"004B",x"A009",x"004C",x"A00A",x"42A1",x"4324",x"42BB",x"004C",x"A00A",x"004D",x"A00A",x"42C2", -- 0620-062F 
  x"A008",x"9004",x"0001",x"004C",x"42EF",x"8FF0",x"004C",x"A00A",x"004B",x"A009",x"004C",x"A00A",x"42A1",x"003C",x"42BB",x"9004", -- 0630-063F 
  x"004C",x"A00A",x"004D",x"A009",x"004C",x"A00A",x"42A1",x"4324",x"42BB",x"A00B",x"004C",x"A00A",x"004D",x"A00A",x"42C2",x"A008", -- 0640-064F 
  x"9004",x"0001",x"004C",x"42EF",x"8FE5",x"004B",x"A00A",x"004C",x"A00A",x"B502",x"42B4",x"B501",x"9003",x"0001",x"004C",x"42EF", -- 0650-065F 
  x"42FA",x"B300",x"A003",x"FFBA",x"E2DE",x"0002",x"47BD",x"430D",x"B502",x"4324",x"42B4",x"9007",x"42FA",x"B300",x"B300",x"B300", -- 0660-066F 
  x"B300",x"0000",x"8023",x"42FA",x"B300",x"B412",x"0000",x"B603",x"42B4",x"9016",x"430D",x"430D",x"B502",x"42A1",x"B502",x"42A1", -- 0670-067F 
  x"42B4",x"9004",x"B300",x"B300",x"0000",x"0000",x"B501",x"9004",x"42AD",x"B412",x"42AD",x"B412",x"42FA",x"42FA",x"42AD",x"8FE7", -- 0680-068F 
  x"B200",x"B300",x"9002",x"FFFF",x"8001",x"0000",x"A003",x"FFCC",x"E2E1",x"0004",x"47BD",x"430D",x"430D",x"0000",x"0051",x"A00A", -- 0690-069F 
  x"0041",x"A00A",x"9003",x"B501",x"A00A",x"A007",x"B501",x"42AD",x"B501",x"A00A",x"B412",x"42AD",x"A00A",x"42FA",x"42FA",x"B603", -- 06A0-06AF 
  x"430D",x"430D",x"4667",x"9003",x"B412",x"A00D",x"B412",x"B502",x"A00D",x"B502",x"A00A",x"A00D",x"A00B",x"A008",x"B502",x"B501", -- 06B0-06BF 
  x"A00A",x"A007",x"0051",x"A00A",x"42BB",x"A00B",x"A008",x"9004",x"B501",x"A00A",x"A007",x"8FDA",x"42FA",x"B300",x"42FA",x"B434", -- 06C0-06CF 
  x"A00D",x"9004",x"B300",x"B300",x"0000",x"0000",x"A003",x"FFC0",x"E2E6",x"0004",x"47BD",x"B412",x"0003",x"A007",x"B412",x"A003", -- 06D0-06DF 
  x"FFF7",x"E2EB",x"0008",x"47BD",x"407F",x"4000",x"A007",x"432D",x"A003",x"FFF7",x"E2F4",x"0006",x"47BD",x"4416",x"004F",x"A00A", -- 06E0-06EF 
  x"0051",x"A00A",x"B502",x"42B4",x"432D",x"0051",x"A009",x"0020",x"4621",x"41E6",x"0001",x"0041",x"A009",x"A003",x"FFEB",x"E2FB", -- 06F0-06FF 
  x"0009",x"47BD",x"004A",x"A00A",x"430D",x"004B",x"A00A",x"430D",x"004C",x"A00A",x"430D",x"004D",x"A00A",x"430D",x"B502",x"A007", -- 0700-070F 
  x"004D",x"A009",x"B501",x"004A",x"A009",x"B501",x"004B",x"A009",x"004C",x"A009",x"0020",x"4621",x"B501",x"901F",x"B603",x"469B", -- 0710-071F 
  x"B501",x"9009",x"430D",x"430D",x"B200",x"42FA",x"42FA",x"46DB",x"B300",x"4338",x"8011",x"B200",x"B603",x"45A4",x"9005",x"B200", -- 0720-072F 
  x"B300",x"0003",x"43F2",x"8008",x"B434",x"B300",x"B412",x"B300",x"0050",x"A00A",x"9001",x"4089",x"8FDD",x"B200",x"42FA",x"004D", -- 0730-073F 
  x"A009",x"42FA",x"004C",x"A009",x"42FA",x"004B",x"A009",x"42FA",x"004A",x"A009",x"A003",x"FFB3",x"E305",x"0004",x"47BD",x"0042", -- 0740-074F 
  x"A00A",x"D002",x"A009",x"0040",x"A00A",x"9006",x"003C",x"4346",x"E30A",x"0004",x"421F",x"8003",x"E30F",x"0002",x"421F",x"439D", -- 0750-075F 
  x"0049",x"A00A",x"0100",x"450F",x"B502",x"A00A",x"003C",x"42BB",x"9002",x"B200",x"802B",x"0040",x"A00A",x"900C",x"003C",x"4346", -- 0760-076F 
  x"E312",x"0003",x"421F",x"4702",x"003C",x"4346",x"E316",x"0004",x"421F",x"801C",x"001B",x"4346",x"005B",x"4346",x"0033",x"4346", -- 0770-077F 
  x"0036",x"4346",x"006D",x"4346",x"4702",x"0050",x"A00A",x"A00D",x"9003",x"E31B",x"0002",x"421F",x"001B",x"4346",x"005B",x"4346", -- 0780-078F 
  x"0033",x"4346",x"0039",x"4346",x"006D",x"4346",x"8FC8",x"A003",x"FFB3",x"E31E",x"0005",x"47BD",x"E324",x"000B",x"421F",x"439D", -- 0790-079F 
  x"439D",x"474F",x"A003",x"FFF5",x"E330",x"0006",x"47BD",x"0000",x"0041",x"A009",x"A003",x"FFF8",x"E337",x"000C",x"47BD",x"42FA", -- 07A0-07AF 
  x"430D",x"A003",x"FFF9",x"E344",x"000A",x"47BD",x"42FA",x"46E4",x"A003",x"FFF9",x"E34F",x"0003",x"47BD",x"42FA",x"0050",x"A00A", -- 07B0-07BF 
  x"9002",x"46E4",x"8001",x"430D",x"A003",x"FFF4",x"E353",x"000A",x"47BD",x"46ED",x"0001",x"0050",x"A009",x"47AE",x"A003",x"FFF6", -- 07C0-07CF 
  x"E35E",x"0008",x"47BD",x"46ED",x"0001",x"0050",x"A009",x"47B5",x"A003",x"FFF6",x"E367",x"0001",x"47BD",x"46ED",x"0001",x"0050", -- 07D0-07DF 
  x"A009",x"47BC",x"A003",x"FFF6",x"E369",x"0001",x"47AF",x"0000",x"0050",x"A009",x"441F",x"407F",x"A003",x"432D",x"47A7",x"A003", -- 07E0-07EF 
  x"FFF3",x"E36B",x"0005",x"47BD",x"4225",x"A003",x"FFFA",x"E371",x"0003",x"47BD",x"47F4",x"A00A",x"9005",x"434D",x"B300",x"434D", -- 07F0-07FF 
  x"B300",x"8006",x"434D",x"4357",x"4346",x"434D",x"4357",x"4346",x"434D",x"4357",x"4346",x"434D",x"4357",x"4346",x"B300",x"A003", -- 0800-080F 
  x"FFE6",x"E375",x"0003",x"47BD",x"E379",x"0001",x"421F",x"0022",x"4346",x"47FA",x"0022",x"4346",x"E37B",x"0001",x"421F",x"A003", -- 0810-081F 
  x"FFF0",x"E37D",x"0005",x"47BD",x"47F4",x"A009",x"0040",x"A00A",x"430D",x"0000",x"0040",x"A009",x"E383",x"0008",x"4219",x"4702", -- 0820-082F 
  x"407F",x"4000",x"A007",x"0010",x"A009",x"439D",x"003C",x"4346",x"E38C",x"0006",x"421F",x"439D",x"E393",x"0002",x"421F",x"0000", -- 0830-083F 
  x"B603",x"A007",x"B501",x"0043",x"42BB",x"9002",x"B300",x"0044",x"A00A",x"4814",x"42AD",x"B501",x"0010",x"42BB",x"9FF1",x"B300", -- 0840-084F 
  x"E396",x"0004",x"421F",x"B501",x"4376",x"E39B",x"0001",x"421F",x"B501",x"000F",x"A007",x"4390",x"0010",x"A007",x"B603",x"42D4", -- 0850-085F 
  x"A00B",x"9FD9",x"B200",x"439D",x"003C",x"4346",x"E39D",x"0007",x"421F",x"42FA",x"0040",x"A009",x"A003",x"FFB3",x"E3A5",x"0005", -- 0860-086F 
  x"4098",x"2F00",x"FFFB",x"E3AB",x"0008",x"47BD",x"2F00",x"A00A",x"B501",x"40A3",x"B501",x"42AD",x"2F00",x"A009",x"A009",x"A003", -- 0870-087F 
  x"FFF2",x"E3B4",x"0004",x"47BD",x"B501",x"900D",x"430D",x"B502",x"A00A",x"B502",x"A009",x"B412",x"42AD",x"B412",x"42AD",x"42FA", -- 0880-088F 
  x"0001",x"42B4",x"8FF1",x"B300",x"B200",x"A003",x"FFEA",x"E3B9",x"0004",x"47BD",x"B434",x"B434",x"B501",x"9009",x"430D",x"B603", -- 0890-089F 
  x"A009",x"0001",x"A007",x"42FA",x"0001",x"42B4",x"8FF5",x"B300",x"B200",x"A003",x"FFEC",x"E3BE",x"0004",x"47BD",x"B412",x"B501", -- 08A0-08AF 
  x"A00A",x"4390",x"0001",x"A007",x"B412",x"0001",x"42B4",x"B501",x"A00D",x"9FF4",x"B300",x"A003",x"FFEE",x"E3C3",x"0003",x"47BD", -- 08B0-08BF 
  x"B603",x"42C2",x"9001",x"B412",x"B300",x"A003",x"FFF6",x"E3C7",x"0003",x"47BD",x"B603",x"42D4",x"9001",x"B412",x"B300",x"A003", -- 08C0-08CF 
  x"FFF6",x"E3CB",x"0003",x"47BD",x"B501",x"A00F",x"9001",x"A000",x"A003",x"FFF7",x"E3CF",x"0006",x"4138",x"A017",x"A003",x"FFFA", -- 08D0-08DF 
  x"E3D6",x"0007",x"4138",x"A018",x"A003",x"FFFA",x"E3DE",x"0009",x"47BD",x"430D",x"A017",x"A018",x"9FFD",x"42FA",x"B300",x"A003", -- 08E0-08EF 
  x"FFF5",x"E3E8",x"0001",x"4098",x"1401",x"FFFB",x"E3EA",x"0001",x"4098",x"1601",x"FFFB",x"E3EC",x"0001",x"4098",x"1801",x"FFFB", -- 08F0-08FF 
  x"E3EE",x"0004",x"47BD",x"0007",x"442C",x"4486",x"A009",x"447D",x"A009",x"4474",x"A009",x"446B",x"A009",x"4462",x"A009",x"445A", -- 0900-090F 
  x"A009",x"4453",x"A009",x"4453",x"A00A",x"446B",x"A00A",x"9001",x"A00B",x"445A",x"A00A",x"4474",x"A00A",x"A007",x"42AD",x"4486", -- 0910-091F 
  x"A00A",x"B502",x"0000",x"489A",x"4486",x"A00A",x"B501",x"4462",x"A00A",x"445A",x"A00A",x"0000",x"B60C",x"A00A",x"B434",x"B434", -- 0920-092F 
  x"447D",x"A00A",x"4474",x"A00A",x"48E9",x"B300",x"A009",x"B300",x"B434",x"0001",x"A007",x"B434",x"0001",x"A007",x"B434",x"FFFF", -- 0930-093F 
  x"A007",x"B501",x"A00D",x"9FE7",x"B300",x"B200",x"4443",x"A003",x"FFB7",x"E3F3",x"0006",x"47BD",x"0007",x"442C",x"4486",x"A009", -- 0940-094F 
  x"447D",x"A009",x"4474",x"A009",x"446B",x"A009",x"4462",x"A009",x"445A",x"A009",x"4453",x"A009",x"4453",x"A00A",x"445A",x"A00A", -- 0950-095F 
  x"4474",x"A00A",x"48C0",x"42AD",x"4486",x"A00A",x"4453",x"A00A",x"446B",x"A00A",x"42BB",x"903C",x"0000",x"445A",x"A00A",x"4474", -- 0960-096F 
  x"A00A",x"48C0",x"0000",x"B434",x"B502",x"B501",x"445A",x"A00A",x"42C2",x"9009",x"4462",x"A00A",x"B501",x"A00A",x"B412",x"42AD", -- 0970-097F 
  x"4462",x"A009",x"8001",x"0000",x"B412",x"4474",x"A00A",x"42C2",x"9009",x"447D",x"A00A",x"B501",x"A00A",x"B412",x"42AD",x"447D", -- 0980-098F 
  x"A009",x"8001",x"0000",x"A001",x"4486",x"A00A",x"B501",x"42AD",x"4486",x"A009",x"A009",x"B434",x"B434",x"0001",x"A007",x"B603", -- 0990-099F 
  x"42B4",x"A00D",x"9FD0",x"B200",x"4486",x"A00A",x"A009",x"8065",x"B412",x"0001",x"42B4",x"B412",x"0001",x"445A",x"A00A",x"4474", -- 09A0-09AF 
  x"A00A",x"48C0",x"0000",x"B434",x"B502",x"B501",x"445A",x"A00A",x"42C2",x"9009",x"4462",x"A00A",x"B501",x"A00A",x"B412",x"42AD", -- 09B0-09BF 
  x"4462",x"A009",x"8001",x"0000",x"B412",x"4474",x"A00A",x"42C2",x"900A",x"447D",x"A00A",x"B501",x"A00A",x"B412",x"42AD",x"447D", -- 09C0-09CF 
  x"A009",x"A00B",x"8001",x"FFFF",x"A001",x"4486",x"A00A",x"B501",x"42AD",x"4486",x"A009",x"A009",x"B434",x"B434",x"0001",x"A007", -- 09D0-09DF 
  x"B603",x"42B4",x"A00D",x"9FCF",x"B200",x"A00D",x"9026",x"B501",x"4486",x"A009",x"B434",x"A00B",x"B434",x"B434",x"0001",x"445A", -- 09E0-09EF 
  x"A00A",x"4474",x"A00A",x"48C0",x"0000",x"B434",x"0000",x"4486",x"A00A",x"A00A",x"A00B",x"A001",x"4486",x"A00A",x"B501",x"42AD", -- 09F0-09FF 
  x"4486",x"A009",x"A009",x"B434",x"B434",x"0001",x"A007",x"B603",x"42B4",x"A00D",x"9FEA",x"B200",x"B300",x"4443",x"A003",x"FF39", -- 0A00-0A0F 
  x"E3FA",x"0004",x"4138",x"A014",x"A003",x"FFFA",x"E3FF",x"0005",x"47BD",x"0010",x"430D",x"A014",x"42FA",x"0001",x"42B4",x"B501", -- 0A10-0A1F 
  x"A00D",x"9FF8",x"B200",x"A003",x"FFF1",x"E405",x"0004",x"47BD",x"0000",x"B434",x"B434",x"4A19",x"A003",x"FFF7",x"E40A",x"0004", -- 0A20-0A2F 
  x"47BD",x"B502",x"A00F",x"9012",x"B412",x"A000",x"B412",x"B501",x"A00F",x"9006",x"A000",x"4A28",x"B412",x"A000",x"B412",x"8005", -- 0A30-0A3F 
  x"4A28",x"A000",x"B412",x"A000",x"B412",x"8008",x"B501",x"A00F",x"9004",x"A000",x"4A28",x"A000",x"8001",x"4A28",x"A003",x"FFDE", -- 0A40-0A4F 
  x"E40F",x"0001",x"47BD",x"4A31",x"B412",x"B300",x"A003",x"FFF8",x"E411",x"0003",x"47BD",x"4A31",x"B300",x"A003",x"FFF9",x"E415", -- 0A50-0A5F 
  x"0004",x"47BD",x"0007",x"442C",x"4486",x"A009",x"447D",x"A009",x"4474",x"A009",x"446B",x"A009",x"4462",x"A009",x"445A",x"A009", -- 0A60-0A6F 
  x"4453",x"A009",x"445A",x"A00A",x"4474",x"A00A",x"42C2",x"900A",x"4453",x"A00A",x"445A",x"A00A",x"4462",x"A00A",x"0000",x"0000", -- 0A70-0A7F 
  x"0000",x"80E1",x"445A",x"A00A",x"0000",x"4462",x"A00A",x"B502",x"A007",x"A00A",x"A00B",x"B502",x"4486",x"A00A",x"A007",x"A009", -- 0A80-0A8F 
  x"0001",x"A007",x"B603",x"42B4",x"A00D",x"9FEF",x"B200",x"4486",x"A00A",x"445A",x"A00A",x"A007",x"4474",x"A00A",x"42B4",x"4462", -- 0A90-0A9F 
  x"A009",x"FFFF",x"4486",x"A00A",x"445A",x"A00A",x"A007",x"A009",x"0001",x"445A",x"42EF",x"445A",x"A00A",x"4474",x"A00A",x"42B4", -- 0AA0-0AAF 
  x"0000",x"4462",x"A00A",x"4474",x"A00A",x"A007",x"A00A",x"A00B",x"4462",x"A00A",x"4474",x"A00A",x"A007",x"0001",x"42B4",x"A00A", -- 0AB0-0ABF 
  x"A00B",x"447D",x"A00A",x"4474",x"A00A",x"A007",x"0001",x"42B4",x"A00A",x"4A19",x"B412",x"B300",x"B501",x"4462",x"A00A",x"4474", -- 0AC0-0ACF 
  x"A00A",x"A007",x"42AD",x"A009",x"0000",x"4462",x"A00A",x"447D",x"A00A",x"4474",x"A00A",x"48E9",x"B200",x"B412",x"B300",x"0000", -- 0AD0-0ADF 
  x"4462",x"A00A",x"4474",x"A00A",x"A007",x"A00A",x"A001",x"4462",x"A00A",x"4474",x"A00A",x"A007",x"A009",x"902C",x"0001",x"4474", -- 0AE0-0AEF 
  x"A00A",x"0000",x"B434",x"B502",x"4462",x"A00A",x"B502",x"A007",x"A00A",x"B412",x"447D",x"A00A",x"A007",x"A00A",x"A00B",x"A001", -- 0AF0-0AFF 
  x"B412",x"430D",x"B502",x"4462",x"A00A",x"A007",x"A009",x"42FA",x"B434",x"B434",x"0001",x"A007",x"B603",x"42B4",x"A00D",x"9FE2", -- 0B00-0B0F 
  x"B200",x"FFFF",x"4462",x"A00A",x"4474",x"A00A",x"A007",x"42AD",x"42EF",x"8FD3",x"FFFF",x"4462",x"42EF",x"0001",x"A007",x"B603", -- 0B10-0B1F 
  x"42B4",x"A00D",x"9F8E",x"B200",x"4474",x"A00A",x"0000",x"4486",x"A00A",x"B502",x"A007",x"A00A",x"A00B",x"B502",x"4486",x"A00A", -- 0B20-0B2F 
  x"A007",x"A009",x"0001",x"A007",x"B603",x"42B4",x"A00D",x"9FEF",x"B200",x"4474",x"A00A",x"4486",x"A00A",x"0001",x"42B4",x"A009", -- 0B30-0B3F 
  x"445A",x"A00A",x"4474",x"A00A",x"42B4",x"4486",x"A00A",x"4474",x"A00A",x"A007",x"A009",x"4453",x"A00A",x"4474",x"A00A",x"4486", -- 0B40-0B4F 
  x"A00A",x"4453",x"A00A",x"446B",x"A00A",x"9001",x"A00B",x"445A",x"A00A",x"4474",x"A00A",x"42B4",x"4486",x"A00A",x"4474",x"A00A", -- 0B50-0B5F 
  x"A007",x"0001",x"A007",x"4443",x"A003",x"FEF9",x"E41A",x"0008",x"4098",x"2F01",x"FFFB",x"E423",x"0008",x"4098",x"2F02",x"FFFB", -- 0B60-0B6F 
  x"E42C",x"0008",x"4098",x"2F03",x"FFFB",x"E435",x"000E",x"4098",x"2F04",x"FFFB",x"E444",x"000C",x"4098",x"2F05",x"FFFB",x"E451", -- 0B70-0B7F 
  x"0006",x"4098",x"2F06",x"FFFB",x"E458",x"000D",x"47BD",x"B502",x"A00D",x"9004",x"B200",x"B300",x"0000",x"8031",x"B603",x"A007", -- 0B80-0B8F 
  x"0001",x"42B4",x"B501",x"A00A",x"A00D",x"A00B",x"9FF9",x"0001",x"A007",x"B502",x"48C0",x"B603",x"42BB",x"9004",x"B200",x"B200", -- 0B90-0B9F 
  x"0000",x"801D",x"B502",x"42B4",x"B502",x"A00A",x"C000",x"A008",x"A00D",x"B502",x"0001",x"42BB",x"A008",x"9003",x"B300",x"A00A", -- 0BA0-0BAF 
  x"8009",x"B502",x"0001",x"42B4",x"A009",x"0001",x"42B4",x"407F",x"4000",x"A00E",x"B412",x"B300",x"B412",x"9001",x"A000",x"A003", -- 0BB0-0BBF 
  x"FFC3",x"E466",x"000C",x"47BD",x"B501",x"A00A",x"B501",x"A00F",x"9003",x"A000",x"FFFF",x"8001",x"0000",x"B434",x"B434",x"B501", -- 0BC0-0BCF 
  x"407F",x"4000",x"A008",x"9009",x"B412",x"B300",x"3FFF",x"A008",x"B501",x"A00A",x"B412",x"42AD",x"8004",x"B502",x"A009",x"0001", -- 0BD0-0BDF 
  x"B412",x"A003",x"FFDE",x"E473",x"000B",x"47BD",x"2F03",x"A00A",x"B603",x"A009",x"42AD",x"B603",x"A007",x"2F03",x"A009",x"B603", -- 0BE0-0BEF 
  x"B412",x"0000",x"489A",x"B412",x"B300",x"2F03",x"A00A",x"2F05",x"A00A",x"42C2",x"A00B",x"9002",x"0369",x"43F2",x"A003",x"FFE3", -- 0BF0-0BFF 
  x"E47F",x"0010",x"47BD",x"2F02",x"A009",x"2F01",x"A009",x"2F01",x"4BC4",x"B502",x"430D",x"2F02",x"4BC4",x"B502",x"42FA",x"A007", -- 0C00-0C0F 
  x"42AD",x"4BE6",x"A003",x"FFEC",x"E490",x"0002",x"47BD",x"4C03",x"494C",x"4B87",x"A003",x"FFF8",x"E493",x"0002",x"47BD",x"A000", -- 0C10-0C1F 
  x"4C17",x"A003",x"FFF9",x"E496",x"0002",x"47BD",x"4C03",x"4903",x"4B87",x"A003",x"FFF8",x"E499",x"0007",x"47AF",x"0051",x"A00A", -- 0C20-0C2F 
  x"0004",x"A007",x"46E4",x"A003",x"FFF6",x"E4A1",x"0005",x"47BD",x"B501",x"A00D",x"9002",x"0000",x"43F2",x"B501",x"2F01",x"A009", -- 0C30-0C3F 
  x"2F01",x"4BC4",x"B434",x"B300",x"B502",x"A007",x"0001",x"42B4",x"A00A",x"B412",x"0001",x"42D4",x"9018",x"0001",x"B502",x"A00F", -- 0C40-0C4F 
  x"A00B",x"9007",x"B412",x"B501",x"A007",x"B412",x"B501",x"4C17",x"8FF5",x"B412",x"B300",x"B501",x"2F06",x"A009",x"B434",x"B502", -- 0C50-0C5F 
  x"4C26",x"B434",x"B434",x"4C26",x"8004",x"B300",x"0001",x"2F06",x"A009",x"4C03",x"4A62",x"4B87",x"430D",x"4B87",x"42FA",x"2F06", -- 0C60-0C6F 
  x"A00A",x"0001",x"42B4",x"9007",x"B412",x"2F06",x"A00A",x"4C38",x"B412",x"B300",x"B412",x"A003",x"FFB8",x"E4A7",x"0004",x"47BD", -- 0C70-0C7F 
  x"0000",x"430D",x"434D",x"B501",x"9007",x"4357",x"4346",x"42FA",x"B300",x"FFFF",x"430D",x"8001",x"B300",x"434D",x"B501",x"4324", -- 0C80-0C8F 
  x"A00E",x"9007",x"4357",x"4346",x"42FA",x"B300",x"FFFF",x"430D",x"8001",x"B300",x"434D",x"B501",x"4324",x"A00E",x"9003",x"4357", -- 0C90-0C9F 
  x"4346",x"8001",x"B300",x"434D",x"4357",x"4346",x"B300",x"42FA",x"B300",x"A003",x"FFD2",x"E4AC",x"0002",x"47BD",x"2F01",x"A009", -- 0CA0-0CAF 
  x"2F01",x"4BC4",x"B434",x"9003",x"E4AF",x"0001",x"421F",x"B502",x"A007",x"0001",x"42B4",x"B501",x"A00A",x"4C80",x"B412",x"0001", -- 0CB0-0CBF 
  x"42B4",x"B412",x"B502",x"900A",x"0001",x"42B4",x"B501",x"A00A",x"4376",x"B412",x"0001",x"42B4",x"B412",x"8FF4",x"B300",x"B300", -- 0CC0-0CCF 
  x"0020",x"4346",x"A003",x"FFD7",x"E4B1",x"0003",x"47BD",x"B412",x"4CAE",x"4CAE",x"A003",x"FFF8",x"E4B5",x"000B",x"4098",x"2F07", -- 0CD0-0CDF 
  x"FFFB",x"E4C1",x"0009",x"4098",x"2F08",x"FFFB",x"E4CB",x"000D",x"47BD",x"2F03",x"A00A",x"A003",x"FFF9",x"E4D9",x"000D",x"47BD", -- 0CE0-0CEF 
  x"2F03",x"A009",x"A003",x"FFF9",x"E4E7",x"000B",x"47BD",x"2F08",x"A00A",x"2F07",x"A009",x"2F03",x"A00A",x"2F08",x"A009",x"A003", -- 0CF0-0CFF 
  x"FFF3",x"E4F3",x"0004",x"47BD",x"2F04",x"A00A",x"2F03",x"A009",x"4CF7",x"4CF7",x"A003",x"FFF5",x"E4F8",x"0003",x"47BD",x"2F01", -- 0D00-0D0F 
  x"A009",x"2F01",x"4BC4",x"B502",x"2F03",x"A00A",x"42AD",x"B412",x"4884",x"2F03",x"A00A",x"42AD",x"B502",x"42AD",x"2F03",x"42EF", -- 0D10-0D1F 
  x"4B87",x"A003",x"FFE9",x"E4FC",x"0003",x"47BD",x"B412",x"4D0F",x"B412",x"4D0F",x"A003",x"FFF7",x"E500",x"0002",x"47BD",x"4CE9", -- 0D20-0D2F 
  x"B434",x"B434",x"4C38",x"B412",x"B300",x"B412",x"4CF0",x"4D0F",x"A003",x"FFF2",x"E503",x"0004",x"47BD",x"4CE9",x"B434",x"B434", -- 0D30-0D3F 
  x"4C38",x"B300",x"B412",x"4CF0",x"4D0F",x"A003",x"FFF3",x"E508",x"0004",x"47BD",x"4CE9",x"B434",x"B434",x"B501",x"9004",x"B412", -- 0D40-0D4F 
  x"B502",x"4D3D",x"8FFA",x"B300",x"B412",x"4CF0",x"4D0F",x"A003",x"FFEE",x"E50D",x"0003",x"47BD",x"4CE9",x"B434",x"B434",x"B603", -- 0D50-0D5F 
  x"4D4A",x"B434",x"B502",x"4D2F",x"B434",x"B434",x"4D2F",x"B434",x"4CF0",x"4D26",x"A003",x"FFED",x"E511",x"0007",x"47BD",x"4CE9", -- 0D60-0D6F 
  x"B434",x"B434",x"0007",x"442C",x"445A",x"A009",x"4453",x"A009",x"0000",x"445A",x"A00A",x"9063",x"B501",x"4462",x"A009",x"0001", -- 0D70-0D7F 
  x"447D",x"A009",x"FFFF",x"4486",x"A009",x"4453",x"A00A",x"4462",x"A00A",x"A007",x"42A1",x"002B",x"42BB",x"9009",x"4462",x"A00A", -- 0D80-0D8F 
  x"42AD",x"4462",x"A009",x"0000",x"4486",x"A009",x"8016",x"4453",x"A00A",x"4462",x"A00A",x"A007",x"42A1",x"002D",x"42BB",x"900D", -- 0D90-0D9F 
  x"4462",x"A00A",x"42AD",x"4462",x"A009",x"0000",x"4486",x"A009",x"447D",x"A00A",x"A000",x"447D",x"A009",x"4486",x"A00A",x"9FD2", -- 0DA0-0DAF 
  x"4462",x"A00A",x"445A",x"A00A",x"42C2",x"9029",x"4453",x"A00A",x"4462",x"A00A",x"A007",x"42A1",x"B501",x"9015",x"457B",x"A00B", -- 0DB0-0DBF 
  x"9007",x"B300",x"445A",x"A00A",x"A000",x"445A",x"A009",x"800A",x"B412",x"0048",x"A00A",x"4C26",x"4C17",x"4462",x"A00A",x"42AD", -- 0DC0-0DCF 
  x"4462",x"A009",x"8005",x"B300",x"4462",x"A00A",x"445A",x"A009",x"4462",x"A00A",x"445A",x"A00A",x"42C2",x"A00B",x"9FD7",x"447D", -- 0DD0-0DDF 
  x"A00A",x"A00F",x"9001",x"A000",x"4462",x"A00A",x"445A",x"A00A",x"42B4",x"B501",x"9006",x"B300",x"4453",x"A00A",x"4462",x"A00A", -- 0DE0-0DEF 
  x"A007",x"4443",x"B434",x"4CF0",x"B412",x"4D0F",x"B412",x"A003",x"FF73",x"E519",x"0002",x"0022",x"41FE",x"4D6F",x"B300",x"A003", -- 0DF0-0DFF 
  x"FFF8",x"E51C",x"0002",x"47BD",x"4CE9",x"B434",x"B434",x"0004",x"442C",x"B501",x"A00F",x"9002",x"0012",x"43F2",x"0002",x"446B", -- 0E00-0E0F 
  x"A009",x"4462",x"A009",x"445A",x"A009",x"0001",x"4462",x"A00A",x"446B",x"A00A",x"4A31",x"4462",x"A009",x"9003",x"445A",x"A00A", -- 0E10-0E1F 
  x"4C26",x"4462",x"A00A",x"9008",x"445A",x"A00A",x"445A",x"A00A",x"4C26",x"445A",x"A009",x"8FEA",x"4443",x"B412",x"4CF0",x"4D0F", -- 0E20-0E2F 
  x"A003",x"FFCF",x"E51F",x"0002",x"47BD",x"0048",x"A00A",x"0010",x"42BB",x"9002",x"4CAE",x"802C",x"4CE9",x"B412",x"B501",x"A00F", -- 0E30-0E3F 
  x"9004",x"A000",x"E522",x"0001",x"421F",x"B501",x"A00D",x"9005",x"E524",x"0002",x"421F",x"B300",x"801A",x"FFFF",x"B412",x"B501", -- 0E40-0E4F 
  x"9004",x"0048",x"A00A",x"4C38",x"8FFA",x"B300",x"B501",x"A00F",x"A00B",x"900A",x"0030",x"A007",x"B501",x"0039",x"42D4",x"9002", -- 0E50-0E5F 
  x"0007",x"A007",x"4346",x"8FF2",x"0020",x"4346",x"B300",x"4CF0",x"A003",x"FFC8",x"E527",x"0003",x"47BD",x"B412",x"4E35",x"4E35", -- 0E60-0E6F 
  x"A003",x"FFF8",x"E52B",x"0006",x"47BD",x"3FFF",x"A008",x"B501",x"42AD",x"B412",x"A00A",x"A003",x"FFF5",x"E532",x"0004",x"47BD", -- 0E70-0E7F 
  x"48D4",x"B501",x"407F",x"4000",x"42C2",x"9003",x"B300",x"0000",x"800A",x"4E75",x"B412",x"B300",x"407F",x"4000",x"42C2",x"9002", -- 0E80-0E8F 
  x"0000",x"8001",x"FFFF",x"A003",x"FFE8",x"E537",x"0001",x"47BD",x"B502",x"4E80",x"9011",x"B412",x"4E75",x"3FFF",x"A008",x"B434", -- 0E90-0E9F 
  x"B603",x"42D4",x"9005",x"B412",x"B300",x"A007",x"A00A",x"8003",x"B200",x"B300",x"0000",x"8003",x"9002",x"B300",x"0000",x"A003", -- 0EA0-0EAF 
  x"FFE4",x"E539",x"0001",x"47BD",x"B603",x"4E98",x"A003",x"FFF9",x"E53B",x"0001",x"47BD",x"B501",x"430D",x"B434",x"B434",x"B502", -- 0EB0-0EBF 
  x"4E80",x"A00D",x"B502",x"A00D",x"A008",x"42FA",x"4E80",x"A00D",x"A008",x"9002",x"B200",x"806F",x"B502",x"4E80",x"A00D",x"9017", -- 0EC0-0ECF 
  x"B501",x"42AD",x"4BE6",x"B434",x"B502",x"A009",x"407F",x"4000",x"B502",x"0001",x"42B4",x"42EF",x"B501",x"430D",x"A007",x"A009", -- 0ED0-0EDF 
  x"42FA",x"0001",x"42B4",x"407F",x"4000",x"A007",x"8054",x"B502",x"4E75",x"3FFF",x"A008",x"B434",x"B603",x"42D4",x"9008",x"B412", -- 0EE0-0EEF 
  x"B300",x"B434",x"430D",x"A007",x"A009",x"42FA",x"801B",x"B501",x"42AD",x"4BE6",x"B412",x"430D",x"B501",x"430D",x"B412",x"4884", -- 0EF0-0EFF 
  x"B300",x"42FA",x"407F",x"4000",x"B502",x"0001",x"42B4",x"42EF",x"B412",x"B502",x"42FA",x"A007",x"A009",x"0001",x"42B4",x"407F", -- 0F00-0F0F 
  x"4000",x"A007",x"4E75",x"3FFF",x"A008",x"B603",x"A007",x"0001",x"42B4",x"A00A",x"A00D",x"B502",x"0001",x"42D4",x"A008",x"9003", -- 0F10-0F1F 
  x"0001",x"42B4",x"8FF2",x"B502",x"A00A",x"4E80",x"A00D",x"B502",x"0001",x"42BB",x"A008",x"9003",x"B300",x"A00A",x"800C",x"B412", -- 0F20-0F2F 
  x"0001",x"42B4",x"B412",x"407F",x"4000",x"A007",x"B502",x"A009",x"407F",x"4000",x"A007",x"A003",x"FF7B",x"E53D",x"0002",x"47BD", -- 0F30-0F3F 
  x"B501",x"4E80",x"9017",x"E540",x"0002",x"421F",x"4E75",x"3FFF",x"A008",x"B502",x"A007",x"B412",x"B603",x"42D4",x"9006",x"B501", -- 0F40-0F4F 
  x"A00A",x"4F40",x"0001",x"A007",x"8FF7",x"B200",x"E543",x"0002",x"421F",x"8001",x"4E35",x"A003",x"FFE0",x"E546",x"0006",x"4098", -- 0F50-0F5F 
  x"2F09",x"FFFB",x"E54D",x"0001",x"47BD",x"2F09",x"A00A",x"D001",x"A00A",x"2F09",x"A009",x"A003",x"FFF5",x"E54F",x"0001",x"47BD", -- 0F60-0F6F 
  x"0000",x"D001",x"A00A",x"0001",x"42B4",x"2F09",x"A00A",x"42B4",x"900A",x"D001",x"A00A",x"0002",x"42B4",x"2F09",x"A00A",x"42B4", -- 0F70-0F7F 
  x"B434",x"4EBB",x"8FEE",x"B412",x"2F09",x"A009",x"A003",x"FFE5",x"E551",x"000B",x"47BD",x"0008",x"442C",x"445A",x"A009",x"4453", -- 0F80-0F8F 
  x"A009",x"0000",x"447D",x"A009",x"0000",x"4486",x"A009",x"4453",x"A00A",x"0001",x"445A",x"A00A",x"4462",x"A009",x"FFFF",x"4462", -- 0F90-0F9F 
  x"42EF",x"448F",x"A009",x"4453",x"A00A",x"4462",x"A00A",x"4E98",x"4462",x"A00A",x"4E98",x"445A",x"A00A",x"446B",x"A009",x"FFFF", -- 0FA0-0FAF 
  x"446B",x"42EF",x"B502",x"446B",x"A00A",x"4E98",x"4462",x"A00A",x"4E98",x"447D",x"A00A",x"446B",x"A00A",x"B434",x"4EBB",x"447D", -- 0FB0-0FBF 
  x"A009",x"B502",x"4462",x"A00A",x"4E98",x"446B",x"A00A",x"4E98",x"4486",x"A00A",x"446B",x"A00A",x"B434",x"4EBB",x"4486",x"A009", -- 0FC0-0FCF 
  x"446B",x"A00A",x"A00D",x"9FDB",x"447D",x"A00A",x"4462",x"A00A",x"4E98",x"448F",x"A00A",x"4C17",x"447D",x"A00A",x"4462",x"A00A", -- 0FD0-0FDF 
  x"B434",x"4EBB",x"447D",x"A009",x"4486",x"A00A",x"4462",x"A00A",x"4E98",x"448F",x"A00A",x"4C1F",x"4486",x"A00A",x"4462",x"A00A", -- 0FE0-0FEF 
  x"B434",x"4EBB",x"4486",x"A009",x"445A",x"A00A",x"446B",x"A009",x"FFFF",x"446B",x"42EF",x"B502",x"446B",x"A00A",x"4E98",x"445A", -- 0FF0-0FFF 
  x"A00A",x"4474",x"A009",x"FFFF",x"4474",x"42EF",x"4CE9",x"B434",x"B434",x"B412",x"B502",x"4474",x"A00A",x"4E98",x"B502",x"4C26", -- 1000-100F 
  x"447D",x"A00A",x"446B",x"A00A",x"4E98",x"4486",x"A00A",x"4474",x"A00A",x"4E98",x"4C26",x"4C1F",x"448F",x"A00A",x"4D2F",x"B43C", -- 1010-101F 
  x"B412",x"4CF0",x"B412",x"4D0F",x"B412",x"4474",x"A00A",x"B434",x"4EBB",x"4474",x"A00A",x"A00D",x"9FD6",x"B434",x"446B",x"A00A", -- 1020-102F 
  x"B434",x"4EBB",x"B412",x"446B",x"A00A",x"A00D",x"9FC1",x"4462",x"A00A",x"A00D",x"9F63",x"4443",x"A003",x"FF4A",x"E55D",x"0005", -- 1030-103F 
  x"47BD",x"0051",x"A00A",x"B501",x"42AD",x"A00A",x"B502",x"0002",x"A007",x"A00A",x"4365",x"0020",x"4346",x"B501",x"A00A",x"9004", -- 1040-104F 
  x"B501",x"A00A",x"A007",x"8FEF",x"B300",x"A003",x"FFE7",x"E563",x"0005",x"47BD",x"0051",x"A00A",x"B501",x"4390",x"B501",x"42AD", -- 1050-105F 
  x"A00A",x"B502",x"0002",x"A007",x"A00A",x"4365",x"0020",x"4346",x"B501",x"A00A",x"9004",x"B501",x"A00A",x"A007",x"8FED",x"B300", -- 1060-106F 
  x"A003",x"FFE5",x"E569",x"0006",x"4098",x"A003",x"FFFB",x"E570",x"0008",x"47BD",x"4416",x"0020",x"4621",x"469B",x"B501",x"9012", -- 1070-107F 
  x"46DB",x"B300",x"42AD",x"4225",x"B412",x"004F",x"A009",x"B501",x"46E4",x"407F",x"A003",x"432D",x"004F",x"A009",x"0001",x"0050", -- 1080-108F 
  x"A009",x"8003",x"B200",x"0003",x"43F2",x"A003",x"FFE0",x"E579",x"0006",x"47BD",x"0020",x"4621",x"469B",x"900E",x"004F",x"A009", -- 1090-109F 
  x"4225",x"B501",x"A00A",x"A007",x"0051",x"A009",x"4225",x"42AD",x"A00A",x"0053",x"A009",x"8004",x"B300",x"E580",x"000F",x"421F", -- 10A0-10AF 
  x"A003",x"FFE5",x"E590",x"000A",x"47BD",x"439D",x"B501",x"0000",x"42BB",x"9003",x"E59B",x"0013",x"421F",x"B501",x"0003",x"42BB", -- 10B0-10BF 
  x"9003",x"E5AF",x"0014",x"421F",x"B501",x"0006",x"42BB",x"9003",x"E5C4",x"0014",x"421F",x"B501",x"0009",x"42BB",x"9003",x"E5D9", -- 10C0-10CF 
  x"0030",x"421F",x"B501",x"0012",x"42BB",x"9003",x"E60A",x"0012",x"421F",x"B501",x"0369",x"42BB",x"9003",x"E61D",x"0013",x"421F", -- 10D0-10DF 
  x"B501",x"1234",x"42BB",x"9003",x"E631",x"004C",x"421F",x"A003",x"FFC9",x"E67E",x"0005",x"47BD",x"47DD",x"4225",x"0003",x"42B4", -- 10E0-10EF 
  x"B501",x"4390",x"A00A",x"42AD",x"B501",x"4390",x"A00A",x"B501",x"4390",x"0040",x"42B4",x"4225",x"B412",x"0007",x"A008",x"0018", -- 10F0-10FF 
  x"A007",x"A009",x"A003",x"FFE5",x"E684",x"0002",x"47BD",x"0007",x"4346",x"E687",x"0008",x"421F",x"A003",x"FFF6",x"E690",x"0002", -- 1100-110F 
  x"47BD",x"0007",x"4346",x"E693",x"0004",x"421F",x"474F",x"A003",x"FFF5",x"E698",x"0002",x"47BD",x"E69B",x"0029",x"421F",x"439D", -- 1110-111F 
  x"FA00",x"0100",x"450F",x"4702",x"E6C5",x"0002",x"421F",x"A003",x"FFF0",x"E6C8",x"0005",x"47BD",x"0049",x"A00A",x"0100",x"450F", -- 1120-112F 
  x"A003",x"FFF7",x"E6CE",x"0007",x"47AF",x"003C",x"4346",x"E6D6",x"0004",x"421F",x"439D",x"512C",x"E6DB",x"0007",x"4219",x"4667", -- 1130-113F 
  x"9FF9",x"003C",x"4346",x"E6E3",x"0003",x"421F",x"A003",x"FFEA",x"E6E7",x"0003",x"47BD",x"0010",x"0048",x"A009",x"A003",x"FFF8", -- 1140-114F 
  x"E6EB",x"0007",x"47BD",x"000A",x"0048",x"A009",x"A003",x"FFF8",x"E6F3",x"0005",x"47BD",x"B501",x"3FFF",x"42D4",x"B502",x"C000", -- 1150-115F 
  x"42C2",x"A00E",x"9002",x"1234",x"43F2",x"432D",x"A003",x"515B",x"A003",x"4D6F",x"A003",x"FFEC",x"E6F9",x"0002",x"47BD",x"4390", -- 1160-116F 
  x"A003",x"FFFA",x"E6FC",x"0002",x"47BD",x"A007",x"A003",x"FFFA",x"E6FF",x"0002",x"47BD",x"42B4",x"A003",x"FFFA",x"E702",x"0002", -- 1170-117F 
  x"47BD",x"42DB",x"A003",x"FFFA",x"E705",x"0002",x"47BD",x"4A53",x"A003",x"FFFA",x"E708",x"0005",x"47BD",x"4A31",x"A003",x"FFFA", -- 1180-118F 
  x"E70E",x"0004",x"47BD",x"4A5B",x"A003",x"FFFA",x"E713",x"0001",x"47BD",x"4F40",x"A003",x"FFFA",x"E715",x"0001",x"47BD",x"4C17", -- 1190-119F 
  x"A003",x"FFFA",x"E717",x"0001",x"47BD",x"4C1F",x"A003",x"FFFA",x"E719",x"0001",x"47BD",x"4C26",x"A003",x"FFFA",x"E71B",x"0001", -- 11A0-11AF 
  x"47BD",x"4D2F",x"A003",x"FFFA",x"E71D",x"0004",x"47BD",x"4C38",x"47DD",x"47DD",x"4A5B",x"4D3D",x"A003",x"FFF6",x"E722",x"0003", -- 11B0-11BF 
  x"47BD",x"4D4A",x"A003",x"FFFA",x"E726",x"0002",x"47BD",x"4D5C",x"A003",x"FFFA",x"E729",x"0001",x"47BD",x"4E04",x"A003",x"FFFA", -- 11C0-11CF 
  x"E72B",x"0001",x"47BD",x"A00A",x"5199",x"A003",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 11D0-11DF 
  others=>x"0000");

-- Textspeicher E000H-FFFFH
type ByteRAMTYPE is array(0 to 8*1024-1) of STD_LOGIC_VECTOR (7 downto 0);
signal ByteRAM: ByteRAMTYPE:=(
  x"28",x"20",x"7B",x"20",x"7D",x"20",x"43",x"4F",x"4D",x"50",x"49",x"4C",x"45",x"20",x"28",x"4C", -- E000-E00F 
  x"49",x"54",x"2C",x"29",x"20",x"4C",x"49",x"54",x"2C",x"20",x"28",x"43",x"4F",x"4E",x"53",x"54", -- E010-E01F 
  x"41",x"4E",x"54",x"3A",x"29",x"20",x"43",x"4F",x"4E",x"53",x"54",x"41",x"4E",x"54",x"20",x"53", -- E020-E02F 
  x"50",x"20",x"52",x"50",x"20",x"50",x"43",x"20",x"58",x"42",x"49",x"54",x"20",x"53",x"4D",x"55", -- E030-E03F 
  x"44",x"47",x"45",x"42",x"49",x"54",x"20",x"52",x"50",x"30",x"20",x"49",x"52",x"41",x"4D",x"41", -- E040-E04F 
  x"44",x"52",x"20",x"4A",x"52",x"41",x"4D",x"41",x"44",x"52",x"20",x"58",x"4F",x"46",x"46",x"20", -- E050-E05F 
  x"43",x"52",x"42",x"5A",x"45",x"49",x"47",x"20",x"43",x"52",x"44",x"50",x"20",x"42",x"41",x"53", -- E060-E06F 
  x"45",x"20",x"54",x"49",x"42",x"20",x"49",x"4E",x"31",x"20",x"49",x"4E",x"32",x"20",x"49",x"4E", -- E070-E07F 
  x"33",x"20",x"49",x"4E",x"34",x"20",x"45",x"52",x"52",x"4F",x"52",x"4E",x"52",x"20",x"44",x"50", -- E080-E08F 
  x"20",x"53",x"54",x"41",x"54",x"20",x"4C",x"46",x"41",x"20",x"42",x"41",x"4E",x"46",x"20",x"42", -- E090-E09F 
  x"5A",x"45",x"49",x"47",x"20",x"44",x"50",x"4D",x"45",x"52",x"4B",x"20",x"43",x"53",x"50",x"20", -- E0A0-E0AF 
  x"4C",x"4F",x"43",x"41",x"4C",x"41",x"44",x"44",x"52",x"20",x"56",x"45",x"52",x"53",x"49",x"4F", -- E0B0-E0BF 
  x"4E",x"20",x"52",x"45",x"54",x"55",x"52",x"4E",x"20",x"28",x"4D",x"43",x"4F",x"44",x"45",x"3A", -- E0C0-E0CF 
  x"29",x"20",x"4D",x"43",x"4F",x"44",x"45",x"20",x"4D",x"49",x"4E",x"55",x"53",x"20",x"55",x"2B", -- E0D0-E0DF 
  x"20",x"55",x"2A",x"20",x"30",x"3D",x"20",x"30",x"4C",x"54",x"20",x"45",x"4D",x"49",x"54",x"43", -- E0E0-E0EF 
  x"4F",x"44",x"45",x"20",x"4E",x"4F",x"54",x"20",x"41",x"4E",x"44",x"20",x"4F",x"52",x"20",x"4B", -- E0F0-E0FF 
  x"45",x"59",x"43",x"4F",x"44",x"45",x"20",x"2B",x"20",x"21",x"20",x"40",x"20",x"53",x"57",x"41", -- E100-E10F 
  x"50",x"20",x"4F",x"56",x"45",x"52",x"20",x"44",x"55",x"50",x"20",x"52",x"4F",x"54",x"20",x"44", -- E110-E11F 
  x"52",x"4F",x"50",x"20",x"32",x"53",x"57",x"41",x"50",x"20",x"32",x"4F",x"56",x"45",x"52",x"20", -- E120-E12F 
  x"32",x"44",x"55",x"50",x"20",x"32",x"44",x"52",x"4F",x"50",x"20",x"4E",x"4F",x"4F",x"50",x"20", -- E130-E13F 
  x"42",x"2C",x"20",x"5A",x"2C",x"20",x"28",x"57",x"4F",x"52",x"44",x"3A",x"29",x"20",x"57",x"4F", -- E140-E14F 
  x"52",x"44",x"3A",x"20",x"22",x"20",x"2E",x"22",x"20",x"48",x"45",x"52",x"45",x"20",x"4A",x"52", -- E150-E15F 
  x"42",x"49",x"54",x"20",x"4A",x"52",x"30",x"42",x"49",x"54",x"20",x"58",x"53",x"45",x"54",x"42", -- E160-E16F 
  x"54",x"20",x"41",x"4C",x"4C",x"4F",x"54",x"20",x"42",x"52",x"41",x"4E",x"43",x"48",x"2C",x"20", -- E170-E17F 
  x"30",x"42",x"52",x"41",x"4E",x"43",x"48",x"2C",x"20",x"42",x"45",x"47",x"49",x"4E",x"20",x"41", -- E180-E18F 
  x"47",x"41",x"49",x"4E",x"20",x"55",x"4E",x"54",x"49",x"4C",x"20",x"49",x"46",x"20",x"45",x"4E", -- E190-E19F 
  x"44",x"5F",x"49",x"46",x"20",x"45",x"4C",x"53",x"45",x"20",x"57",x"48",x"49",x"4C",x"45",x"20", -- E1A0-E1AF 
  x"52",x"45",x"50",x"45",x"41",x"54",x"20",x"43",x"40",x"20",x"43",x"21",x"20",x"31",x"2B",x"20", -- E1B0-E1BF 
  x"2D",x"20",x"3D",x"20",x"4C",x"54",x"20",x"3E",x"20",x"2A",x"20",x"42",x"59",x"45",x"20",x"42", -- E1C0-E1CF 
  x"59",x"45",x"20",x"20",x"2B",x"21",x"20",x"52",x"3E",x"20",x"3E",x"52",x"20",x"52",x"20",x"2C", -- E1D0-E1DF 
  x"20",x"45",x"58",x"45",x"43",x"55",x"54",x"45",x"20",x"4B",x"45",x"59",x"20",x"45",x"4D",x"49", -- E1E0-E1EF 
  x"54",x"20",x"53",x"48",x"4C",x"31",x"36",x"20",x"44",x"49",x"47",x"20",x"54",x"59",x"50",x"45", -- E1F0-E1FF 
  x"20",x"48",x"47",x"2E",x"20",x"48",x"2E",x"20",x"2E",x"20",x"3F",x"20",x"43",x"52",x"20",x"66", -- E200-E20F 
  x"6C",x"3E",x"20",x"2F",x"66",x"6C",x"3E",x"20",x"66",x"72",x"3E",x"20",x"2F",x"66",x"72",x"3E", -- E210-E21F 
  x"20",x"46",x"45",x"48",x"4C",x"45",x"52",x"54",x"45",x"58",x"54",x"20",x"44",x"49",x"53",x"41", -- E220-E22F 
  x"42",x"4C",x"45",x"20",x"77",x"65",x"69",x"74",x"65",x"72",x"20",x"6E",x"61",x"63",x"68",x"20", -- E230-E23F 
  x"54",x"61",x"73",x"74",x"65",x"20",x"45",x"53",x"43",x"41",x"50",x"45",x"20",x"20",x"45",x"52", -- E240-E24F 
  x"52",x"4F",x"52",x"20",x"3F",x"3F",x"3F",x"20",x"46",x"45",x"48",x"4C",x"45",x"52",x"54",x"45", -- E250-E25F 
  x"58",x"54",x"20",x"45",x"52",x"52",x"4F",x"52",x"20",x"2D",x"20",x"46",x"65",x"68",x"6C",x"65", -- E260-E26F 
  x"72",x"20",x"4E",x"75",x"6D",x"6D",x"65",x"72",x"20",x"20",x"43",x"53",x"50",x"21",x"20",x"43", -- E270-E27F 
  x"53",x"50",x"3F",x"20",x"4C",x"4F",x"43",x"41",x"4C",x"20",x"45",x"4E",x"44",x"5F",x"4C",x"4F", -- E280-E28F 
  x"43",x"41",x"4C",x"20",x"4C",x"30",x"20",x"4C",x"31",x"20",x"4C",x"32",x"20",x"4C",x"33",x"20", -- E290-E29F 
  x"4C",x"34",x"20",x"4C",x"35",x"20",x"4C",x"36",x"20",x"4C",x"37",x"20",x"27",x"20",x"49",x"4E", -- E2A0-E2AF 
  x"43",x"52",x"34",x"20",x"4B",x"45",x"59",x"5F",x"49",x"4E",x"54",x"20",x"4B",x"45",x"59",x"43", -- E2B0-E2BF 
  x"4F",x"44",x"45",x"32",x"20",x"45",x"58",x"50",x"45",x"43",x"54",x"20",x"44",x"49",x"47",x"49", -- E2C0-E2CF 
  x"54",x"20",x"4E",x"55",x"4D",x"42",x"45",x"52",x"20",x"57",x"4F",x"52",x"44",x"20",x"5A",x"3D", -- E2D0-E2DF 
  x"20",x"46",x"49",x"4E",x"44",x"20",x"4C",x"43",x"46",x"41",x"20",x"43",x"4F",x"4D",x"50",x"49", -- E2E0-E2EF 
  x"4C",x"45",x"2C",x"20",x"43",x"52",x"45",x"41",x"54",x"45",x"20",x"49",x"4E",x"54",x"45",x"52", -- E2F0-E2FF 
  x"50",x"52",x"45",x"54",x"20",x"51",x"55",x"49",x"54",x"20",x"2F",x"6F",x"6B",x"3E",x"20",x"6F", -- E300-E30F 
  x"6B",x"20",x"6F",x"6B",x"3E",x"20",x"2F",x"6F",x"6B",x"3E",x"20",x"6F",x"6B",x"20",x"53",x"54", -- E310-E31F 
  x"41",x"52",x"54",x"20",x"46",x"4F",x"52",x"54",x"59",x"2D",x"46",x"4F",x"52",x"54",x"48",x"20", -- E320-E32F 
  x"53",x"4D",x"55",x"44",x"47",x"45",x"20",x"28",x"49",x"4D",x"4D",x"45",x"44",x"49",x"41",x"54", -- E330-E33F 
  x"45",x"3A",x"29",x"20",x"28",x"43",x"4F",x"4D",x"50",x"49",x"4C",x"45",x"3A",x"29",x"20",x"28", -- E340-E34F 
  x"3A",x"29",x"20",x"49",x"4D",x"4D",x"45",x"44",x"49",x"41",x"54",x"45",x"3A",x"20",x"43",x"4F", -- E350-E35F 
  x"4D",x"50",x"49",x"4C",x"45",x"3A",x"20",x"3A",x"20",x"3B",x"20",x"44",x"55",x"42",x"49",x"54", -- E360-E36F 
  x"20",x"4C",x"47",x"2E",x"20",x"4E",x"47",x"2E",x"20",x"78",x"20",x"2C",x"20",x"44",x"55",x"4D", -- E370-E37F 
  x"50",x"5A",x"20",x"27",x"20",x"53",x"54",x"41",x"52",x"54",x"20",x"20",x"44",x"55",x"4D",x"50", -- E380-E38F 
  x"5A",x"3E",x"20",x"20",x"20",x"20",x"20",x"2D",x"2D",x"20",x"20",x"2D",x"20",x"2F",x"44",x"55", -- E390-E39F 
  x"4D",x"50",x"5A",x"3E",x"20",x"52",x"41",x"4D",x"50",x"31",x"20",x"56",x"41",x"52",x"49",x"41", -- E3A0-E3AF 
  x"42",x"4C",x"45",x"20",x"4D",x"4F",x"56",x"45",x"20",x"46",x"49",x"4C",x"4C",x"20",x"44",x"55", -- E3B0-E3BF 
  x"4D",x"50",x"20",x"4D",x"41",x"58",x"20",x"4D",x"49",x"4E",x"20",x"41",x"42",x"53",x"20",x"4D", -- E3C0-E3CF 
  x"55",x"4C",x"54",x"5F",x"49",x"20",x"4D",x"55",x"4C",x"54",x"5F",x"49",x"49",x"20",x"53",x"55", -- E3D0-E3DF 
  x"50",x"45",x"52",x"4D",x"55",x"4C",x"54",x"20",x"41",x"20",x"42",x"20",x"43",x"20",x"53",x"4D", -- E3E0-E3EF 
  x"55",x"4C",x"20",x"41",x"44",x"44",x"49",x"45",x"52",x"20",x"44",x"49",x"33",x"32",x"20",x"44", -- E3F0-E3FF 
  x"49",x"56",x"33",x"32",x"20",x"2F",x"4D",x"4F",x"44",x"20",x"2F",x"4D",x"4F",x"44",x"20",x"2F", -- E400-E40F 
  x"20",x"4D",x"4F",x"44",x"20",x"53",x"44",x"49",x"56",x"20",x"4F",x"50",x"45",x"52",x"41",x"4E", -- E410-E41F 
  x"44",x"31",x"20",x"4F",x"50",x"45",x"52",x"41",x"4E",x"44",x"32",x"20",x"45",x"52",x"47",x"45", -- E420-E42F 
  x"42",x"4E",x"49",x"53",x"20",x"5A",x"41",x"48",x"4C",x"45",x"4E",x"53",x"50",x"45",x"49",x"43", -- E430-E43F 
  x"48",x"45",x"52",x"20",x"53",x"50",x"45",x"49",x"43",x"48",x"45",x"52",x"45",x"4E",x"44",x"45", -- E440-E44F 
  x"20",x"53",x"43",x"48",x"49",x"45",x"42",x"20",x"53",x"4C",x"58",x"2D",x"3E",x"45",x"52",x"47", -- E450-E45F 
  x"45",x"42",x"4E",x"49",x"53",x"20",x"4F",x"50",x"45",x"52",x"41",x"4E",x"44",x"2D",x"3E",x"53", -- E460-E46F 
  x"4C",x"58",x"20",x"53",x"50",x"45",x"49",x"43",x"48",x"45",x"52",x"48",x"4F",x"4C",x"20",x"32", -- E470-E47F 
  x"4F",x"50",x"45",x"52",x"41",x"4E",x"44",x"45",x"4E",x"2D",x"3E",x"32",x"53",x"4C",x"58",x"20", -- E480-E48F 
  x"4E",x"2B",x"20",x"4E",x"2D",x"20",x"4E",x"2A",x"20",x"52",x"45",x"43",x"55",x"52",x"53",x"45", -- E490-E49F 
  x"20",x"4E",x"2F",x"4D",x"4F",x"44",x"20",x"48",x"47",x"30",x"2E",x"20",x"4E",x"2E",x"20",x"2D", -- E4A0-E4AF 
  x"20",x"4E",x"42",x"2E",x"20",x"42",x"4C",x"4F",x"43",x"4B",x"41",x"4E",x"46",x"41",x"4E",x"47", -- E4B0-E4BF 
  x"20",x"42",x"4C",x"4F",x"43",x"4B",x"45",x"4E",x"44",x"45",x"20",x"4E",x"45",x"42",x"45",x"4E", -- E4C0-E4CF 
  x"52",x"45",x"43",x"48",x"4E",x"55",x"4E",x"47",x"20",x"48",x"41",x"55",x"50",x"54",x"52",x"45", -- E4D0-E4DF 
  x"43",x"48",x"4E",x"55",x"4E",x"47",x"20",x"52",x"45",x"43",x"48",x"45",x"4E",x"42",x"4C",x"4F", -- E4E0-E4EF 
  x"43",x"4B",x"20",x"49",x"4E",x"49",x"54",x"20",x"41",x"2B",x"30",x"20",x"42",x"2B",x"30",x"20", -- E4F0-E4FF 
  x"4E",x"2F",x"20",x"4E",x"4D",x"4F",x"44",x"20",x"4E",x"47",x"47",x"54",x"20",x"4E",x"42",x"4B", -- E500-E50F 
  x"20",x"4E",x"4E",x"55",x"4D",x"42",x"45",x"52",x"20",x"4E",x"22",x"20",x"4E",x"5E",x"20",x"4E", -- E510-E51F 
  x"2E",x"20",x"2D",x"20",x"30",x"20",x"20",x"4E",x"42",x"2E",x"20",x"5A",x"45",x"52",x"4C",x"45", -- E520-E52F 
  x"47",x"20",x"4F",x"42",x"4A",x"3F",x"20",x"4C",x"20",x"47",x"20",x"48",x"20",x"4F",x"2E",x"20", -- E530-E53F 
  x"5B",x"20",x"20",x"5D",x"20",x"20",x"53",x"50",x"4D",x"45",x"52",x"4B",x"20",x"5B",x"20",x"5D", -- E540-E54F 
  x"20",x"49",x"4E",x"56",x"45",x"52",x"54",x"49",x"45",x"52",x"45",x"4E",x"20",x"56",x"4C",x"49", -- E550-E55F 
  x"53",x"54",x"20",x"57",x"4C",x"49",x"53",x"54",x"20",x"52",x"45",x"54",x"55",x"52",x"4E",x"20", -- E560-E56F 
  x"52",x"45",x"50",x"4C",x"41",x"43",x"45",x"3A",x"20",x"46",x"4F",x"52",x"47",x"45",x"54",x"20", -- E570-E57F 
  x"6E",x"69",x"63",x"68",x"74",x"20",x"67",x"65",x"66",x"75",x"6E",x"64",x"65",x"6E",x"20",x"20", -- E580-E58F 
  x"46",x"45",x"48",x"4C",x"45",x"52",x"54",x"45",x"58",x"54",x"20",x"44",x"69",x"76",x"69",x"73", -- E590-E59F 
  x"69",x"6F",x"6E",x"20",x"64",x"75",x"72",x"63",x"68",x"20",x"4E",x"75",x"6C",x"6C",x"20",x"57", -- E5A0-E5AF 
  x"6F",x"72",x"74",x"20",x"6E",x"69",x"63",x"68",x"74",x"20",x"64",x"65",x"66",x"69",x"6E",x"69", -- E5B0-E5BF 
  x"65",x"72",x"74",x"20",x"45",x"69",x"6E",x"67",x"61",x"62",x"65",x"7A",x"65",x"69",x"6C",x"65", -- E5C0-E5CF 
  x"20",x"7A",x"75",x"20",x"6C",x"61",x"6E",x"67",x"20",x"53",x"74",x"72",x"75",x"6B",x"74",x"75", -- E5D0-E5DF 
  x"72",x"66",x"65",x"68",x"6C",x"65",x"72",x"20",x"69",x"6E",x"20",x"49",x"46",x"20",x"45",x"4E", -- E5E0-E5EF 
  x"44",x"5F",x"49",x"46",x"20",x"42",x"45",x"47",x"49",x"4E",x"20",x"55",x"4E",x"54",x"49",x"4C", -- E5F0-E5FF 
  x"20",x"44",x"4F",x"20",x"4C",x"4F",x"4F",x"50",x"20",x"20",x"6E",x"65",x"67",x"61",x"74",x"69", -- E600-E60F 
  x"76",x"65",x"72",x"20",x"45",x"78",x"70",x"6F",x"6E",x"65",x"6E",x"74",x"20",x"5A",x"61",x"68", -- E610-E61F 
  x"6C",x"65",x"6E",x"73",x"70",x"65",x"69",x"63",x"68",x"65",x"72",x"20",x"76",x"6F",x"6C",x"6C", -- E620-E62F 
  x"20",x"67",x"72",x"6F",x"C3",x"9F",x"65",x"20",x"67",x"61",x"6E",x"7A",x"65",x"20",x"5A",x"61", -- E630-E63F 
  x"68",x"6C",x"65",x"6E",x"20",x"6B",x"6F",x"6D",x"70",x"69",x"6C",x"69",x"65",x"72",x"65",x"6E", -- E640-E64F 
  x"20",x"67",x"65",x"68",x"74",x"20",x"6D",x"6F",x"6D",x"65",x"6E",x"74",x"61",x"6E",x"20",x"6E", -- E650-E65F 
  x"69",x"63",x"68",x"74",x"2C",x"20",x"73",x"69",x"65",x"68",x"65",x"20",x"54",x"45",x"53",x"54", -- E660-E66F 
  x"46",x"55",x"45",x"52",x"4E",x"45",x"55",x"45",x"53",x"2E",x"54",x"58",x"54",x"20",x"53",x"54", -- E670-E67F 
  x"52",x"47",x"3A",x"20",x"5E",x"47",x"20",x"2F",x"31",x"78",x"50",x"49",x"45",x"50",x"2F",x"20", -- E680-E68F 
  x"5E",x"46",x"20",x"51",x"55",x"49",x"54",x"20",x"5E",x"41",x"20",x"41",x"6E",x"67",x"65",x"68", -- E690-E69F 
  x"61",x"6C",x"74",x"65",x"6E",x"20",x"66",x"C3",x"BC",x"72",x"20",x"67",x"65",x"6E",x"61",x"75", -- E6A0-E6AF 
  x"20",x"65",x"69",x"6E",x"65",x"20",x"45",x"69",x"6E",x"67",x"61",x"62",x"65",x"7A",x"65",x"69", -- E6B0-E6BF 
  x"6C",x"65",x"3A",x"20",x"20",x"6F",x"6B",x"20",x"51",x"55",x"45",x"52",x"59",x"20",x"28",x"2A", -- E6C0-E6CF 
  x"52",x"45",x"4D",x"2A",x"29",x"20",x"2F",x"6F",x"6B",x"3E",x"20",x"28",x"2A",x"45",x"4E",x"44", -- E6D0-E6DF 
  x"2A",x"29",x"20",x"6F",x"6B",x"3E",x"20",x"48",x"45",x"58",x"20",x"44",x"45",x"43",x"49",x"4D", -- E6E0-E6EF 
  x"41",x"4C",x"20",x"4E",x"4C",x"49",x"54",x"2C",x"20",x"4D",x"2E",x"20",x"4D",x"2B",x"20",x"4D", -- E6F0-E6FF 
  x"2D",x"20",x"4D",x"2A",x"20",x"4D",x"2F",x"20",x"4D",x"2F",x"4D",x"4F",x"44",x"20",x"4D",x"4D", -- E700-E70F 
  x"4F",x"44",x"20",x"2E",x"20",x"2B",x"20",x"2D",x"20",x"2A",x"20",x"2F",x"20",x"2F",x"4D",x"4F", -- E710-E71F 
  x"44",x"20",x"47",x"47",x"54",x"20",x"42",x"4B",x"20",x"5E",x"20",x"3F",x"20",x"00",x"00",x"00", -- E720-E72F 
  others=>x"00");

-- Daten 2C00H-2FFFH
type VarRAMTYPE is array(0 to 1024-1) of STD_LOGIC_VECTOR (15 downto 0);
shared variable VarRAM: VarRAMTYPE:=(
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C00-2C0F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C10-2C1F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C20-2C2F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C30-2C3F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C40-2C4F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C50-2C5F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C60-2C6F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C70-2C7F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C80-2C8F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C90-2C9F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2CA0-2CAF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2CB0-2CBF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2CC0-2CCF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2CD0-2CDF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2CE0-2CEF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2CF0-2CFF 
  x"0000",x"0000",x"0000",x"0000",x"0055",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D00-2D0F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D10-2D1F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D20-2D2F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D30-2D3F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D40-2D4F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D50-2D5F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D60-2D6F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D70-2D7F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D80-2D8F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D90-2D9F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2DA0-2DAF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2DB0-2DBF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2DC0-2DCF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2DD0-2DDF 
  x"FFCE",x"012C",x"FF38",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2DE0-2DEF 
  x"0032",x"FED4",x"0190",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2DF0-2DFF 
  x"000F",x"FFC4",x"0032",x"FFC4",x"0140",x"FED4",x"0032",x"FED4",x"012C",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E00-2E0F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E10-2E1F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E20-2E2F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E30-2E3F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E40-2E4F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E50-2E5F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E60-2E6F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E70-2E7F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E80-2E8F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E90-2E9F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2EA0-2EAF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2EB0-2EBF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2EC0-2ECF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2ED0-2EDF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2EE0-2EEF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2EF0-2EFF 
  x"2F0A",x"0000",x"0000",x"140C",x"1400",x"2000",x"0001",x"1400",x"1400",x"0000",x"0000",x"2EE0",x"0000",x"0000",x"0000",x"0000", -- 2F00-2F0F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F10-2F1F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F20-2F2F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F30-2F3F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F40-2F4F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F50-2F5F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F60-2F6F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F70-2F7F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F80-2F8F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F90-2F9F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2FA0-2FAF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2FB0-2FBF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2FC0-2FCF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0301",x"0301",x"0301",x"0301",x"0301",x"0301",x"0301",x"0301", -- 2FD0-2FDF 
  x"0301",x"0301",x"0301",x"0301",x"0446",x"0446",x"0000",x"0001",x"0301",x"0083",x"02C9",x"0301",x"0301",x"068E",x"0301",x"0083", -- 2FE0-2FEF 
  x"0301",x"0301",x"0301",x"0083",x"0348",x"036F",x"0220",x"02BC",x"0845",x"FFFF",x"072A",x"FB05",x"FB06",x"FB00",x"FB00",x"0774", -- 2FF0-2FFF 
  others=>x"0000");

-- Rueckkehrstapel 3FC0-3FFFH, TRUE_DUAL_PORT
type RetRAMTYPE is array(0 to 63) of STD_LOGIC_VECTOR (15 downto 0);
shared variable RetRAM: RetRAMTYPE:=(
  others=>x"0000");

-- diese Funktion übernimmt von SP nur die beiden niedrigsten Bits
  function P(SP : integer) return integer is begin
--    return CONV_INTEGER(CONV_UNSIGNED(SP,2));
    return SP mod 4;
    end;

-- alles Signale um die Stapel-RAM's zu machen.
signal HOLE_VOM_STAPEL,STORE_ZUM_STAPEL,ADRESSE_ZUM_STAPEL: REG;
signal WE_ZUM_STAPEL: STD_LOGIC_VECTOR (3 downto 0);
type STAPELTYPE is array(0 to 31) of STD_LOGIC_VECTOR (15 downto 0);
signal stap1,stap2,stap3,stap0: STAPELTYPE:=(others=>x"0000");
-- Rueckkehrstapel
signal RPC,RPCC: STD_LOGIC_VECTOR (15 downto 0);
signal RP: STD_LOGIC_VECTOR (15 downto 0):=x"4000"; --auch RP0 auf 4000H setzen.
signal RW: STD_LOGIC;
-- kompletten Speicher anschliessen
signal PC_ZUM_ProgRAM,PD_VOM_ProgRAM: STD_LOGIC_VECTOR (15 downto 0);
signal STORE_ZUM_RAM,EXFET,ADRESSE_ZUM_RAM: STD_LOGIC_VECTOR (15 downto 0);
signal FETCH_VOM_ProgRAM,FETCH_VOM_ByteRAM,FETCH_VOM_VarRAM,FETCH_VOM_RetRAM: STD_LOGIC_VECTOR (15 downto 0);
signal WE_ZUM_RAM,WE_ZUM_ProgRAM,WE_ZUM_ByteRAM,WE_ZUM_VarRAM,WE_ZUM_RetRAM: STD_LOGIC;
-- fuer EMIT-Ausgabe
signal EMIT_ABGESCHICKT_LOCAL,EMIT_ANGEKOMMEN_RUHEND,XOFF_INPUT_L: STD_LOGIC:='0';
signal KEY_ANGEKOMMEN_LOCAL,KEY_ABGESCHICKT_RUHEND,KEY_ABGESCHICKT_MERK: STD_LOGIC:='0';
signal KEY_BYTE_RUHEND: STD_LOGIC_VECTOR (7 downto 0);


begin

process begin wait until (CLK_I'event and CLK_I='1'); --ruhende Eingangsdaten für FortyForthprocessor
  EMIT_ANGEKOMMEN_RUHEND<=EMIT_ANGEKOMMEN;
  KEY_BYTE_RUHEND<=KEY_BYTE;
  KEY_ABGESCHICKT_RUHEND<=KEY_ABGESCHICKT;
  end process;
  

process -- FortyForthProcessor
variable PC,PD,ADR,DAT,DIST: STD_LOGIC_VECTOR (15 downto 0):=x"0000";
variable WE: STD_LOGIC;
variable SP: integer:=0;
variable R: REG:=(others=>x"0000");
-- Stapeleintraege benennen
variable A,B,C,D: STD_LOGIC_VECTOR (15 downto 0):=x"0000";
variable T: integer range 0 to 4;
variable W: STD_LOGIC_VECTOR (3 downto 0);
-- fuer Umstapeln 
variable STAK: STD_LOGIC_VECTOR (7 downto 0);
-- fuer Rechenoperationen mit Uebertrag
variable U: STD_LOGIC_VECTOR (31 downto 0);
-- fuer Division
variable UBIT: STD_LOGIC;
-- fuer Supermult
variable SUMME: STD_LOGIC_VECTOR (31 downto 0);

begin wait until (CLK_I'event and CLK_I='0'); PC_SIM<=PC;--Simulation
  -- ob ein KEY aingetroffen ist --
  if KEY_ABGESCHICKT_MERK/=KEY_ABGESCHICKT_RUHEND then 
    KEY_ABGESCHICKT_MERK<=KEY_ABGESCHICKT_RUHEND;
    PD:=x"4026";
    PC:=PC;
    else
      PD:=PD_VOM_ProgRAM;
      PC:=PC+1;
      end if;                                           -- Simulation --
  WE:='0';                                              PD_SIM<=PD;
  DIST:=PD(11)&PD(11)&PD(11)&PD(11)&PD(11 downto 0);    SP_SIM<=SP;
  -- oberste 4 Stapeleintraege entnehmen
  R:=HOLE_VOM_STAPEL;                                   -- Simulation --
  A:=R(P(SP-1));                                        A_SIM<=A;
  B:=R(P(SP-2));                                        B_SIM<=B;
  C:=R(P(SP-3));                                        C_SIM<=C;
  D:=R(P(SP-4));                                        D_SIM<=D;
  T:=0;
  -- Rueckkehrstapel
  RW<='0';
 
  if PD(15 downto 13)="010" then                 -- 4000-5FFF Unterprogrammaufruf
    RPC<=PC;PC:=PD and x"3FFF";RP<=RP-1;RW<='1';
    elsif PD(15 downto 12)=x"8" then PC:=PC+DIST;-- 8000-8FFF relativer Sprung
    elsif PD(15 downto 12)=x"9" then             -- 9000-9FFF bedingter relativer Sprung
      if A=x"0000" then PC:=PC+DIST; end if; SP:=SP-1;
    elsif PD=x"A003" then PC:=RPCC;RP<=RP+1;     -- ; Rückkehr aus Unterprogramm
    elsif PD=x"A00D" then -- 0= Vergleich ob gleich Null
      if A=x"0000" then A:=x"FFFF"; 
        else A:=x"0000"; end if;
      T:=1;
    elsif PD=x"A00F" then -- 0< Vergleich ob kleiner Null
      if A>=x"8000" then A:=x"FFFF";
        else A:=x"0000"; end if;
      T:=1;
    elsif PD=x"A000" then -- MINUS Vorzeichen wechseln
      A:=(not A)+1;
      T:=1;
    elsif PD=x"A00B" then -- NOT Bitweises Komplement
      A:=not A;
      T:=1;
    elsif PD=x"A008" then -- AND Bitweises Und
      A:=B and A; 
      T:=1;
      SP:=SP-1;
    elsif PD=x"A00E" then -- OR Bitweises Oder
      A:=B or A; 
      T:=1;
      SP:=SP-1;
    elsif PD=x"A007" then -- + Addition
      A:=B+A; 
      T:=1;
      SP:=SP-1;
    elsif PD=x"A001" then -- U+ Addition mit Übertrag
      U:=(x"0000"&C)+(x"0000"&B)+(x"0000"&A);
      B:=U(31 downto 16);
      A:=U(15 downto 0);
      T:=2;
      SP:=SP-1;
    elsif PD=x"A002" then -- U* Multiplikation mit Übertrag
      U:=(x"0000"&C)+B*A;
      B:=U(31 downto 16);
      A:=U(15 downto 0);
      T:=2;
      SP:=SP-1;
    elsif PD=x"A005" then -- EMIT Zeichen ausgeben
      if (EMIT_ABGESCHICKT_LOCAL=EMIT_ANGEKOMMEN_RUHEND) and XOFF_INPUT_L='0' then
        EMIT_BYTE<=A(7 downto 0);
        EMIT_ABGESCHICKT_LOCAL<=not EMIT_ANGEKOMMEN_RUHEND;
        T:=0;
        SP:=SP-1;
        else PC:=PC-1; end if; -- warten
    elsif PD=x"A009" then -- STORE Speicheradresse beschreiben
      case A is
        when x"D000" => KEY_ANGEKOMMEN_LOCAL<=not KEY_ANGEKOMMEN_LOCAL;
        when x"D001" => SP:=CONV_INTEGER(B);
        when x"D002" => RP<=B;
        when x"D003" => PC:=B;
        when others => ADR:=A;DAT:=B;WE:='1' ;
        end case;
      T:=0;
      SP:=SP-2;
    elsif PD=x"A00A" then -- FETCH Speicheradresse lesen
      case A is
        when x"D000" => A:=x"00"&KEY_BYTE_RUHEND;
        when x"D001" => A:=CONV_STD_LOGIC_VECTOR(SP-1,16);
        when x"D002" => A:=RP;
        when x"D003" => A:=PC;
        when others => A:=EXFET;
        end case;
      T:=1;
    elsif PD=x"A014" then -- DI32 DIVISION_MIT_REST 32B/16B=16R/16Q
      UBIT:=C(15);
      C:=C(14 downto 0)&B(15);
      B:=B(14 downto 0)&'0';
      if (UBIT&C)>=('0'&A) then
        C:=C-A;
        B(0):='1';
        end if;
      T:=3;
    elsif PD=x"A017" then -- MULT_I
      --     D    C    B    A        RetRAM
      --     c    ü   adr1 adr2      i
      -- c   ü   erg1 adr2 adr1      i-1
      SUMME:=(D*EXFET)+(x"0000"&C);
      C:=A;A:=B;B:=C;
      D:=SUMME(31 downto 16); 
      C:=SUMME(15 downto 0);
      RPC<=RPCC-1; RW<='1';
      T:=4; SP:=SP+1;
    elsif PD=x"A018" then -- MULT_II
      --     D    C     B      A         RetRAM
      -- c   ü1  erg1   adr2   adr1      i-1
      -- c   ü2  adr1+1 adr2+1 i-1       i-1
      SUMME:=(D&C)+(x"0000"&EXFET);
      D:=SUMME(31 downto 16); 
      DAT:=SUMME(15 downto 0);
      ADR:=A;
      WE:='1';
      C:=A+1;
      B:=B+1;
      if RPCC=x"0000" then A:=x"FFFF"; else A:=x"0000"; end if;
      T:=4;
    elsif PD(15 downto 12)=x"B" then           -- B000-BFFF Umstapeln
      STAK:="00000000";
      if PD(7)='1' then STAK:=STAK(5 downto 0)&"11"; T:=T+1; end if;
      if PD(6)='1' then STAK:=STAK(5 downto 0)&"10"; T:=T+1; end if;
      if PD(5)='1' then STAK:=STAK(5 downto 0)&"01"; T:=T+1; end if;
      if PD(4)='1' then STAK:=STAK(5 downto 0)&"00"; T:=T+1; end if;
      if PD(3)='1' then STAK:=STAK(5 downto 0)&"11"; T:=T+1; end if;
      if PD(2)='1' then STAK:=STAK(5 downto 0)&"10"; T:=T+1; end if;
      if PD(1)='1' then STAK:=STAK(5 downto 0)&"01"; T:=T+1; end if;
      if PD(0)='1' then STAK:=STAK(5 downto 0)&"00"; T:=T+1; end if;
      A:=R(P(SP-1-CONV_INTEGER(STAK(1 downto 0))));
      B:=R(P(SP-1-CONV_INTEGER(STAK(3 downto 2))));
      C:=R(P(SP-1-CONV_INTEGER(STAK(5 downto 4))));
      D:=R(P(SP-1-CONV_INTEGER(STAK(7 downto 6))));
      SP:=SP+CONV_INTEGER(PD(11 downto 8))-4;
    else A:=PD; SP:=SP+1; T:=1; end if;                    -- LIT
    
  -- oberste T Stapeleintraege zurückspeichern
  W:="0000";
  if T/=0 then R(P(SP-1)):=A; W(P(SP-1)):='1';
    if T/=1 then R(P(SP-2)):=B; W(P(SP-2)):='1';
      if T/=2 then R(P(SP-3)):=C; W(P(SP-3)):='1';
        if T/=3 then R(P(SP-4)):=D; W(P(SP-4)):='1';
          end if; end if; end if; end if;
  -- Ausgabeadresse zum VarRAMAM zusammenbasteln
  ADRESSE_ZUM_STAPEL(0)<=CONV_STD_LOGIC_VECTOR(SP-1,16);
  ADRESSE_ZUM_STAPEL(1)<=CONV_STD_LOGIC_VECTOR(SP-2,16);
  ADRESSE_ZUM_STAPEL(2)<=CONV_STD_LOGIC_VECTOR(SP-3,16);
  ADRESSE_ZUM_STAPEL(3)<=CONV_STD_LOGIC_VECTOR(SP-4,16);
  STORE_ZUM_STAPEL<=R;
  WE_ZUM_STAPEL<=W;
  -- ADR, DAT, WE, PC
  if WE='1' then ADRESSE_ZUM_RAM<=ADR; else ADRESSE_ZUM_RAM<=R(P(SP-1)); end if;
  STORE_ZUM_RAM<=DAT;
  WE_ZUM_RAM<=WE;
  PC_ZUM_ProgRAM<=PC;
  end process;

ADR_O<=ADRESSE_ZUM_RAM;
DAT_O<=STORE_ZUM_RAM;
WE_O<=WE_ZUM_RAM;
EMIT_ABGESCHICKT<=EMIT_ABGESCHICKT_LOCAL;
KEY_ANGEKOMMEN<=KEY_ANGEKOMMEN_LOCAL;

-- hier werden die Lesedaten der unterschiedlichen Speicher zusammengefuehrt
EXFET<=FETCH_VOM_ProgRAM when ADRESSE_ZUM_RAM(15 downto 13)="000" else
       FETCH_VOM_VarRAM when ADRESSE_ZUM_RAM(15 downto 10)="001011" else
       FETCH_VOM_RetRAM when ADRESSE_ZUM_RAM(15 downto 6)="0011111111" else
       x"00"&FETCH_VOM_ByteRAM(7 downto 0) when ADRESSE_ZUM_RAM(15 downto 13)="111" else
       DAT_I;

-- hier wird WE auf die unterschiedlichen Speicher aufgeteilt
WE_ZUM_ProgRAM<=WE_ZUM_RAM when ADRESSE_ZUM_RAM(15 downto 13)="000" else '0';
WE_ZUM_VarRAM  <=WE_ZUM_RAM when ADRESSE_ZUM_RAM(15 downto 10)="001011" else '0';
WE_ZUM_RetRAM<=WE_ZUM_RAM when ADRESSE_ZUM_RAM(15 downto 6)="0011111111" else '0';
WE_ZUM_ByteRAM<=WE_ZUM_RAM when ADRESSE_ZUM_RAM(15 downto 13)="111" else '0';


process -- Programmspeicher 0000H-1FFFH,
begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_ProgRAM='1' then 
    ProgRAM(CONV_INTEGER(ADRESSE_ZUM_RAM(12 downto 0)))<=STORE_ZUM_RAM; 
    FETCH_VOM_ProgRAM<=STORE_ZUM_RAM; 
	  else
      FETCH_VOM_ProgRAM<=ProgRAM(CONV_INTEGER(ADRESSE_ZUM_RAM(12 downto 0)));
      end if;
  PD_VOM_ProgRAM<=ProgRAM(CONV_INTEGER(PC_ZUM_ProgRAM(12 downto 0)));
  end process;

process -- Textspeicher E000H-FFFFH
begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_ByteRAM='1' then 
    ByteRAM(CONV_INTEGER(ADRESSE_ZUM_RAM(12 downto 0)))<=STORE_ZUM_RAM(7 downto 0); 
    FETCH_VOM_ByteRAM<=STORE_ZUM_RAM; 
	 else
      FETCH_VOM_ByteRAM<=x"00"&ByteRAM(CONV_INTEGER(ADRESSE_ZUM_RAM(12 downto 0)));
      end if;
  end process;

process -- Daten 2C00H-2FFFH
begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_VarRAM='1' then 
    VarRAM(CONV_INTEGER(ADRESSE_ZUM_RAM(9 downto 0))):=STORE_ZUM_RAM; 
    FETCH_VOM_VarRAM<=STORE_ZUM_RAM; 
      else
      FETCH_VOM_VarRAM<=VarRAM(CONV_INTEGER(ADRESSE_ZUM_RAM(9 downto 0)));
      end if;
  FETCH_VOM_VarRAM<=VarRAM(CONV_INTEGER(ADRESSE_ZUM_RAM(9 downto 0)));
  end process;

process --Rueckkehrstapel 3FC0-3FFFH, TRUE_DUAL_PORT
begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_RetRAM='1' then 
    RetRAM(CONV_INTEGER(ADRESSE_ZUM_RAM(5 downto 0))):=STORE_ZUM_RAM; 
    FETCH_VOM_RetRAM<=STORE_ZUM_RAM; 
      else
      FETCH_VOM_RetRAM<=RetRAM(CONV_INTEGER(ADRESSE_ZUM_RAM(5 downto 0)));
      end if;
  FETCH_VOM_RetRAM<=RetRAM(CONV_INTEGER(ADRESSE_ZUM_RAM(5 downto 0)));
  end process;
process begin wait until (CLK_I'event and CLK_I='1');
  if RW='1' then
    RetRAM(CONV_INTEGER(RP(5 downto 0))):=RPC;
    RPCC<=RPC;
     else
      RPCC<=RetRAM(CONV_INTEGER(RP(5 downto 0)));
    end if;
  end process;

--StapelRAM:
process begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_STAPEL(0)='1' then
    stap0(CONV_INTEGER(ADRESSE_ZUM_STAPEL(0)(6 downto 2)))<=STORE_ZUM_STAPEL(0);
    HOLE_VOM_STAPEL(0)<=STORE_ZUM_STAPEL(0);
     else
      HOLE_VOM_STAPEL(0)<=stap0(CONV_INTEGER(ADRESSE_ZUM_STAPEL(0)(6 downto 2)));
    end if;
  end process;
process begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_STAPEL(1)='1' then
    stap1(CONV_INTEGER(ADRESSE_ZUM_STAPEL(1)(6 downto 2)))<=STORE_ZUM_STAPEL(1);
    HOLE_VOM_STAPEL(1)<=STORE_ZUM_STAPEL(1);
     else
      HOLE_VOM_STAPEL(1)<=stap1(CONV_INTEGER(ADRESSE_ZUM_STAPEL(1)(6 downto 2)));
    end if;
  end process;
process begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_STAPEL(2)='1' then
    stap2(CONV_INTEGER(ADRESSE_ZUM_STAPEL(2)(6 downto 2)))<=STORE_ZUM_STAPEL(2);
    HOLE_VOM_STAPEL(2)<=STORE_ZUM_STAPEL(2);
     else
      HOLE_VOM_STAPEL(2)<=stap2(CONV_INTEGER(ADRESSE_ZUM_STAPEL(2)(6 downto 2)));
    end if;
  end process;
process begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_STAPEL(3)='1' then
    stap3(CONV_INTEGER(ADRESSE_ZUM_STAPEL(3)(6 downto 2)))<=STORE_ZUM_STAPEL(3);
    HOLE_VOM_STAPEL(3)<=STORE_ZUM_STAPEL(3);
     else
      HOLE_VOM_STAPEL(3)<=stap3(CONV_INTEGER(ADRESSE_ZUM_STAPEL(3)(6 downto 2)));
    end if;
  end process;

end Step_9;
