library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity FortyForthProcessor is
  Port (
    CLK_I: in STD_LOGIC;
    DAT_I: in STD_LOGIC_VECTOR (15 downto 0);
    ADR_O: out STD_LOGIC_VECTOR (15 downto 0);
    DAT_O: out STD_LOGIC_VECTOR (15 downto 0);
    WE_O: out STD_LOGIC;
    
    -- EMIT --
    EMIT_ABGESCHICKT: out STD_LOGIC;
    EMIT_BYTE: out STD_LOGIC_VECTOR (7 downto 0);
    EMIT_ANGEKOMMEN: in STD_LOGIC;
    
     -- EMIT --
    KEY_ABGESCHICKT: in STD_LOGIC;
    KEY_BYTE: in STD_LOGIC_VECTOR (7 downto 0);
    KEY_ANGEKOMMEN: out STD_LOGIC;

   -- nur zur Simulation und Fehlersuche:
    PC_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    PD_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    SP_SIM: out integer;
    A_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    B_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    C_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    D_SIM: out STD_LOGIC_VECTOR (15 downto 0)
    );
end FortyForthProcessor;

architecture Step_9 of FortyForthProcessor is

constant SHA: STD_LOGIC_VECTOR (10*16-1 downto 0):=
  x"39de37159cb53472ef59b9bdf699180c9c43d52a";
type REG is array(0 to 3) of STD_LOGIC_VECTOR (15 downto 0);
type RAMTYPE is array(0 to 8*1024-1) of STD_LOGIC_VECTOR (15 downto 0);
-- Programmspeicher 0000H-1FFFH
signal ProgRAM: RAMTYPE:=(
  x"4010",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 0000-000F 
  x"4763",x"A003",x"4481",x"A003",x"4000",x"A003",x"4000",x"A003",x"4000",x"A003",x"4000",x"A003",x"4000",x"A003",x"0010",x"A003", -- 0010-001F 
  x"0000",x"3000",x"0001",x"4776",x"0029",x"45E8",x"B200",x"A003",x"FFF8",x"3002",x"0001",x"4776",x"0000",x"2F10",x"A009",x"A003", -- 0020-002F 
  x"FFF8",x"3004",x"0001",x"4784",x"0001",x"2F10",x"A009",x"A003",x"FFF8",x"3006",x"0007",x"4776",x"0020",x"45E8",x"4662",x"46A2", -- 0030-003F 
  x"B300",x"46AB",x"A003",x"FFF5",x"300E",x"0006",x"477D",x"42C6",x"B501",x"4279",x"42D9",x"A00A",x"A003",x"FFF6",x"3015",x"0004", -- 0040-004F 
  x"4784",x"51DB",x"A003",x"42A0",x"B502",x"C000",x"428E",x"A00E",x"9001",x"4046",x"42F9",x"A003",x"FFF1",x"301A",x"000B",x"477D", -- 0050-005F 
  x"42C6",x"A00A",x"2F10",x"A00A",x"9001",x"4051",x"A003",x"FFF5",x"3026",x"0008",x"4784",x"46B4",x"405F",x"42F9",x"476E",x"A003", -- 0060-006F 
  x"FFF7",x"302F",x"0006",x"4060",x"2800",x"FFFB",x"3036",x"0002",x"4060",x"2801",x"FFFB",x"3039",x"0002",x"4060",x"2802",x"FFFB", -- 0070-007F 
  x"303C",x"0002",x"4060",x"2803",x"FFFB",x"303F",x"0004",x"4060",x"2F00",x"FFFB",x"3044",x"0009",x"4060",x"2F01",x"FFFB",x"304E", -- 0080-008F 
  x"0003",x"4060",x"2F02",x"FFFB",x"3052",x"0007",x"4060",x"2F03",x"FFFB",x"305A",x"0007",x"4060",x"2F04",x"FFFB",x"3062",x"0004", -- 0090-009F 
  x"4060",x"2F05",x"FFFB",x"3067",x"0007",x"4060",x"2F06",x"FFFB",x"306F",x"0004",x"4060",x"2F07",x"FFFB",x"3074",x"0004",x"4060", -- 00A0-00AF 
  x"2F08",x"FFFB",x"3079",x"0003",x"4060",x"2F09",x"FFFB",x"307D",x"0003",x"4060",x"2F0A",x"FFFB",x"3081",x"0003",x"4060",x"2F0B", -- 00B0-00BF 
  x"FFFB",x"3085",x"0003",x"4060",x"2F0C",x"FFFB",x"3089",x"0003",x"4060",x"2F0D",x"FFFB",x"308D",x"0007",x"4060",x"2F0E",x"FFFB", -- 00C0-00CF 
  x"3095",x"0002",x"4060",x"2F0F",x"FFFB",x"3098",x"0004",x"4060",x"2F10",x"FFFB",x"309D",x"0003",x"4060",x"2F11",x"FFFB",x"30A1", -- 00D0-00DF 
  x"0004",x"4060",x"2F12",x"FFFB",x"30A6",x"0005",x"4060",x"2F13",x"FFFB",x"30AC",x"0006",x"4060",x"2F14",x"FFFB",x"30B3",x"0003", -- 00E0-00EF 
  x"4060",x"2F15",x"FFFB",x"30B7",x"0005",x"4060",x"2F16",x"FFFB",x"30BD",x"000C",x"4060",x"2F17",x"FFFB",x"30CA",x"0007",x"4060", -- 00F0-00FF 
  x"01BE",x"FFFB",x"30D2",x"0006",x"4060",x"A003",x"FFFB",x"30D9",x"0008",x"477D",x"42C6",x"2F10",x"A00A",x"9003",x"A00A",x"42F9", -- 0100-010F 
  x"8001",x"4304",x"A003",x"FFF3",x"30E2",x"0005",x"4784",x"46B4",x"4109",x"42F9",x"4047",x"A003",x"42F9",x"476E",x"A003",x"FFF4", -- 0110-011F 
  x"30E8",x"0005",x"410A",x"A000",x"A003",x"FFFA",x"30EE",x"0002",x"410A",x"A001",x"A003",x"FFFA",x"30F1",x"0002",x"410A",x"A002", -- 0120-012F 
  x"A003",x"FFFA",x"30F4",x"0002",x"410A",x"A00D",x"A003",x"FFFA",x"30F7",x"0003",x"410A",x"A00F",x"A003",x"FFFA",x"30FB",x"0008", -- 0130-013F 
  x"410A",x"A005",x"A003",x"FFFA",x"3104",x"0003",x"410A",x"A00B",x"A003",x"FFFA",x"3108",x"0003",x"410A",x"A008",x"A003",x"FFFA", -- 0140-014F 
  x"310C",x"0002",x"410A",x"A00E",x"A003",x"FFFA",x"310F",x"0001",x"410A",x"A007",x"A003",x"FFFA",x"3111",x"0001",x"410A",x"A009", -- 0150-015F 
  x"A003",x"FFFA",x"3113",x"0001",x"410A",x"A00A",x"A003",x"FFFA",x"3115",x"0004",x"410A",x"B412",x"A003",x"FFFA",x"311A",x"0004", -- 0160-016F 
  x"410A",x"B502",x"A003",x"FFFA",x"311F",x"0003",x"410A",x"B501",x"A003",x"FFFA",x"3123",x"0003",x"410A",x"B434",x"A003",x"FFFA", -- 0170-017F 
  x"3127",x"0004",x"410A",x"B300",x"A003",x"FFFA",x"312C",x"0005",x"410A",x"B43C",x"A003",x"FFFA",x"3132",x"0005",x"410A",x"B60C", -- 0180-018F 
  x"A003",x"FFFA",x"3138",x"0004",x"410A",x"B603",x"A003",x"FFFA",x"313D",x"0005",x"410A",x"B200",x"A003",x"FFFA",x"3143",x"0004", -- 0190-019F 
  x"410A",x"8000",x"A003",x"FFFA",x"3148",x"0002",x"4784",x"2F13",x"A00A",x"A009",x"0001",x"2F13",x"42BB",x"A003",x"FFF5",x"314B", -- 01A0-01AF 
  x"0002",x"4784",x"2F13",x"A00A",x"4051",x"B501",x"42F9",x"B412",x"B501",x"A00A",x"41A7",x"4279",x"B412",x"0001",x"4280",x"B501", -- 01B0-01BF 
  x"A00D",x"9FF5",x"B200",x"0020",x"41A7",x"A003",x"FFE8",x"314E",x"0007",x"477D",x"45E8",x"2F10",x"A00A",x"9003",x"41B2",x"42C6", -- 01C0-01CF 
  x"46AB",x"A003",x"FFF4",x"3156",x"0005",x"4784",x"46B4",x"0001",x"2F10",x"A009",x"42F9",x"41C9",x"FFFF",x"2F15",x"42BB",x"A003", -- 01D0-01DF 
  x"FFF2",x"315C",x"0001",x"0022",x"41CA",x"A003",x"FFFA",x"315E",x"0002",x"0022",x"41CA",x"4335",x"A003",x"FFF9",x"3161",x"0004", -- 01E0-01EF 
  x"4784",x"2F0F",x"A00A",x"A003",x"FFF9",x"3166",x"0005",x"4784",x"0008",x"A003",x"FFFA",x"316C",x"0006",x"4784",x"0009",x"A003", -- 01F0-01FF 
  x"FFFA",x"3173",x"0006",x"4784",x"1000",x"42A7",x"B412",x"0FFF",x"A008",x"A00E",x"A003",x"FFF5",x"317A",x"0005",x"4784",x"2F0F", -- 0200-020F 
  x"42BB",x"A003",x"FFF9",x"3180",x"0007",x"4784",x"41F1",x"4279",x"4280",x"41F8",x"4204",x"42F9",x"A003",x"FFF5",x"3188",x"0008", -- 0210-021F 
  x"4784",x"41F1",x"4279",x"4280",x"41FE",x"4204",x"42F9",x"A003",x"FFF5",x"3191",x"0005",x"4776",x"41F1",x"A003",x"FFFA",x"3197", -- 0220-022F 
  x"0005",x"4776",x"4216",x"A003",x"FFFA",x"319D",x"0005",x"4776",x"4221",x"A003",x"FFFA",x"31A3",x"0002",x"4776",x"41FE",x"0001", -- 0230-023F 
  x"420F",x"41F1",x"A003",x"FFF7",x"31A6",x"0006",x"4776",x"41F1",x"B502",x"4280",x"B434",x"4204",x"B412",x"0001",x"4280",x"A009", -- 0240-024F 
  x"A003",x"FFF2",x"31AD",x"0004",x"4776",x"0001",x"420F",x"4246",x"41F8",x"41F1",x"A003",x"FFF6",x"31B2",x"0005",x"4776",x"423D", -- 0250-025F 
  x"A003",x"FFFA",x"31B8",x"0006",x"4776",x"B434",x"4231",x"4246",x"A003",x"FFF8",x"31BF",x"0002",x"4784",x"A00A",x"A003",x"FFFA", -- 0260-026F 
  x"31C2",x"0002",x"4784",x"A009",x"A003",x"FFFA",x"31C5",x"0002",x"4784",x"0001",x"A007",x"A003",x"FFF9",x"31C8",x"0001",x"4784", -- 0270-027F 
  x"A000",x"A007",x"A003",x"FFF9",x"31CA",x"0001",x"4784",x"4280",x"A00D",x"A003",x"FFF9",x"31CC",x"0002",x"4784",x"4047",x"8000", -- 0280-028F 
  x"A007",x"B412",x"A00B",x"4047",x"8000",x"A007",x"0000",x"A001",x"B300",x"A00D",x"A00B",x"A003",x"FFEE",x"31CF",x"0001",x"4784", -- 0290-029F 
  x"B412",x"428E",x"A003",x"FFF9",x"31D1",x"0001",x"4784",x"0000",x"B434",x"B434",x"A002",x"B412",x"B300",x"A003",x"FFF5",x"31D3", -- 02A0-02AF 
  x"0003",x"4784",x"31D7",x"0004",x"41EB",x"8FFC",x"A003",x"FFF7",x"31DC",x"0002",x"4784",x"B412",x"B502",x"A00A",x"A007",x"B412", -- 02B0-02BF 
  x"A009",x"A003",x"FFF5",x"31DF",x"0002",x"4784",x"2802",x"A00A",x"4279",x"A00A",x"2802",x"A00A",x"4279",x"2802",x"B603",x"A00A", -- 02C0-02CF 
  x"A00A",x"B412",x"A009",x"A009",x"A003",x"FFED",x"31E2",x"0002",x"4784",x"2802",x"A00A",x"B501",x"FFFF",x"A007",x"2802",x"B603", -- 02D0-02DF 
  x"A00A",x"A00A",x"B412",x"B501",x"FFFF",x"A007",x"2802",x"A009",x"A009",x"A009",x"A009",x"A003",x"FFE9",x"31E5",x"0001",x"4784", -- 02E0-02EF 
  x"2802",x"A00A",x"4279",x"A00A",x"A003",x"FFF7",x"31E7",x"0001",x"4784",x"2F0F",x"A00A",x"A009",x"0001",x"2F0F",x"42BB",x"A003", -- 02F0-02FF 
  x"FFF5",x"31E9",x"0007",x"4784",x"2803",x"A009",x"A003",x"FFF9",x"31F1",x"0003",x"4784",x"8000",x"44B0",x"A00B",x"9002",x"B300", -- 0300-030F 
  x"8FFA",x"A003",x"FFF5",x"31F5",x"0004",x"4784",x"0141",x"4304",x"A003",x"FFF9",x"31FA",x"0005",x"4784",x"0000",x"B412",x"0010", -- 0310-031F 
  x"A002",x"B412",x"A003",x"FFF6",x"3200",x"0003",x"4784",x"B501",x"000A",x"428E",x"9001",x"8002",x"0007",x"A007",x"0030",x"A007", -- 0320-032F 
  x"A003",x"FFF2",x"3204",x"0004",x"4784",x"B501",x"9009",x"B412",x"B501",x"426D",x"4316",x"4279",x"B412",x"0001",x"4280",x"8FF5", -- 0330-033F 
  x"B200",x"A003",x"FFEF",x"3209",x"0003",x"4784",x"431D",x"4327",x"4316",x"431D",x"4327",x"4316",x"431D",x"4327",x"4316",x"431D", -- 0340-034F 
  x"4327",x"4316",x"B300",x"A003",x"FFEE",x"320D",x"0002",x"4784",x"4346",x"0020",x"4316",x"A003",x"FFF8",x"3210",x"0001",x"4784", -- 0350-035F 
  x"4358",x"A003",x"FFFA",x"3212",x"0001",x"4784",x"A00A",x"4360",x"A003",x"FFF9",x"3214",x"0002",x"4784",x"2F07",x"A00A",x"2F0F", -- 0360-036F 
  x"A00A",x"4280",x"2F10",x"A00A",x"A00D",x"A00B",x"A00E",x"2F00",x"A00A",x"A00D",x"A00B",x"A008",x"9028",x"003C",x"4316",x"3217", -- 0370-037F 
  x"0003",x"41EB",x"2F07",x"A00A",x"4360",x"2F06",x"A00A",x"4360",x"003C",x"4316",x"321B",x"0004",x"41EB",x"003C",x"4316",x"3220", -- 0380-038F 
  x"0003",x"41EB",x"2F0F",x"A00A",x"4360",x"2F13",x"A00A",x"4360",x"003C",x"4316",x"3224",x"0004",x"41EB",x"2F0F",x"A00A",x"2F07", -- 0390-039F 
  x"A009",x"2F13",x"A00A",x"2F06",x"A009",x"000A",x"4316",x"A003",x"FFC1",x"3229",x"000A",x"4784",x"A003",x"FFFB",x"3234",x"0007", -- 03A0-03AF 
  x"4784",x"436D",x"323C",x"0019",x"41EB",x"0020",x"4316",x"0008",x"4316",x"430B",x"001B",x"4287",x"9FF8",x"A003",x"FFEF",x"3256", -- 03B0-03BF 
  x"0005",x"4784",x"B501",x"2F0E",x"A009",x"0000",x"2F10",x"A009",x"436D",x"2F0A",x"A00A",x"2F0C",x"A00A",x"2F0A",x"A00A",x"4280", -- 03C0-03CF 
  x"0001",x"4280",x"4335",x"325C",x"0003",x"41EB",x"3260",x"000A",x"41E5",x"46C9",x"436D",x"326B",x"0016",x"41EB",x"4360",x"43B1", -- 03D0-03DF 
  x"4716",x"A003",x"FFDC",x"3282",x"0004",x"4784",x"2801",x"A00A",x"2F15",x"A009",x"A003",x"FFF7",x"3287",x"0004",x"4784",x"2801", -- 03E0-03EF 
  x"A00A",x"2F15",x"A00A",x"4280",x"9002",x"0009",x"43C2",x"A003",x"FFF3",x"328C",x"0005",x"4784",x"0001",x"A007",x"2F17",x"A00A", -- 03F0-03FF 
  x"B502",x"4280",x"B501",x"2F17",x"A009",x"A009",x"A003",x"FFF1",x"3292",x"0009",x"4784",x"2F17",x"A00A",x"B501",x"A00A",x"A007", -- 0400-040F 
  x"2F17",x"A009",x"A003",x"FFF4",x"329C",x"0002",x"4784",x"2F17",x"A00A",x"0001",x"A007",x"A003",x"FFF7",x"329F",x"0002",x"4784", -- 0410-041F 
  x"2F17",x"A00A",x"0002",x"A007",x"A003",x"FFF7",x"32A2",x"0002",x"4784",x"2F17",x"A00A",x"0003",x"A007",x"A003",x"FFF7",x"32A5", -- 0420-042F 
  x"0002",x"4784",x"2F17",x"A00A",x"0004",x"A007",x"A003",x"FFF7",x"32A8",x"0002",x"4784",x"2F17",x"A00A",x"0005",x"A007",x"A003", -- 0430-043F 
  x"FFF7",x"32AB",x"0002",x"4784",x"2F17",x"A00A",x"0006",x"A007",x"A003",x"FFF7",x"32AE",x"0002",x"4784",x"2F17",x"A00A",x"0007", -- 0440-044F 
  x"A007",x"A003",x"FFF7",x"32B1",x"0002",x"4784",x"2F17",x"A00A",x"0008",x"A007",x"A003",x"FFF7",x"32B4",x"0001",x"4776",x"0020", -- 0450-045F 
  x"45E8",x"4662",x"46A2",x"B300",x"4279",x"2F10",x"A00A",x"9001",x"4051",x"A003",x"FFF1",x"32B6",x"0005",x"4784",x"B501",x"A00A", -- 0460-046F 
  x"0001",x"A007",x"B501",x"03FF",x"A008",x"0000",x"4287",x"9002",x"0400",x"4280",x"B412",x"A009",x"A003",x"FFED",x"32BC",x"0007", -- 0470-047F 
  x"4784",x"2800",x"A00A",x"B501",x"0008",x"428E",x"9009",x"0018",x"A007",x"A00A",x"B501",x"9002",x"B501",x"4304",x"B300",x"8018", -- 0480-048F 
  x"2F03",x"A00A",x"A009",x"2F03",x"446E",x"2F03",x"A00A",x"2F04",x"A00A",x"4280",x"03FF",x"A008",x"0080",x"42A0",x"9009",x"2F05", -- 0490-049F 
  x"A00A",x"A00D",x"9005",x"FFFF",x"2F05",x"A009",x"0013",x"4316",x"0000",x"2800",x"A009",x"A003",x"FFD1",x"32C4",x"0008",x"4784", -- 04A0-04AF 
  x"2F04",x"A00A",x"2F03",x"A00A",x"4287",x"9003",x"0000",x"0000",x"8018",x"2F04",x"A00A",x"A00A",x"FFFF",x"2F04",x"446E",x"2F03", -- 04B0-04BF 
  x"A00A",x"2F04",x"A00A",x"4280",x"03FF",x"A008",x"0020",x"428E",x"9008",x"2F05",x"A00A",x"9005",x"0000",x"2F05",x"A009",x"0011", -- 04C0-04CF 
  x"4316",x"A003",x"FFDA",x"32CD",x"0006",x"4784",x"0005",x"43FC",x"4429",x"A009",x"4420",x"A009",x"4420",x"A00A",x"443B",x"A009", -- 04D0-04DF 
  x"430B",x"B501",x"0014",x"4287",x"9004",x"B300",x"4420",x"A00A",x"426D",x"B501",x"007F",x"4287",x"9002",x"B300",x"0008",x"B501", -- 04E0-04EF 
  x"0008",x"4287",x"9012",x"443B",x"A00A",x"4420",x"A00A",x"428E",x"900C",x"FFFF",x"4420",x"42BB",x"0001",x"4429",x"42BB",x"0008", -- 04F0-04FF 
  x"4316",x"0020",x"4316",x"0008",x"4316",x"B501",x"0020",x"428E",x"9001",x"8012",x"FFFF",x"4429",x"42BB",x"4429",x"A00A",x"A00F", -- 0500-050F 
  x"9002",x"0006",x"43C2",x"B501",x"4316",x"B501",x"4420",x"A00A",x"4273",x"0001",x"4420",x"42BB",x"B501",x"0020",x"428E",x"B502", -- 0510-051F 
  x"0008",x"4287",x"A00B",x"A008",x"B412",x"001B",x"4287",x"A00B",x"A008",x"4429",x"A00A",x"A00D",x"A00E",x"9FB2",x"0020",x"4316", -- 0520-052F 
  x"443B",x"A00A",x"4420",x"A00A",x"443B",x"A00A",x"4280",x"B603",x"A007",x"0000",x"B412",x"4273",x"440B",x"A003",x"FF94",x"32D4", -- 0530-053F 
  x"0005",x"4784",x"B501",x"0030",x"428E",x"A00B",x"B502",x"003A",x"428E",x"A008",x"B502",x"0041",x"428E",x"A00B",x"A00E",x"B501", -- 0540-054F 
  x"9015",x"B412",x"0030",x"4280",x"B501",x"000A",x"428E",x"A00B",x"9002",x"0007",x"4280",x"B501",x"2F08",x"A00A",x"428E",x"A00B", -- 0550-055F 
  x"9004",x"B300",x"B300",x"0000",x"0000",x"B412",x"A003",x"FFD7",x"32DA",x"0006",x"4784",x"51DD",x"A003",x"4420",x"A009",x"4417", -- 0560-056F 
  x"A009",x"0000",x"4420",x"A00A",x"9063",x"B501",x"4429",x"A009",x"0001",x"4444",x"A009",x"FFFF",x"444D",x"A009",x"4417",x"A00A", -- 0570-057F 
  x"4429",x"A00A",x"A007",x"426D",x"002B",x"4287",x"9009",x"4429",x"A00A",x"4279",x"4429",x"A009",x"0000",x"444D",x"A009",x"8016", -- 0580-058F 
  x"4417",x"A00A",x"4429",x"A00A",x"A007",x"426D",x"002D",x"4287",x"900D",x"4429",x"A00A",x"4279",x"4429",x"A009",x"0000",x"444D", -- 0590-059F 
  x"A009",x"4444",x"A00A",x"A000",x"4444",x"A009",x"444D",x"A00A",x"9FD2",x"4429",x"A00A",x"4420",x"A00A",x"428E",x"9029",x"4417", -- 05A0-05AF 
  x"A00A",x"4429",x"A00A",x"A007",x"426D",x"B501",x"9015",x"4542",x"A00B",x"9007",x"B300",x"4420",x"A00A",x"A000",x"4420",x"A009", -- 05B0-05BF 
  x"800A",x"B412",x"2F08",x"A00A",x"42A7",x"A007",x"4429",x"A00A",x"4279",x"4429",x"A009",x"8005",x"B300",x"4429",x"A00A",x"4420", -- 05C0-05CF 
  x"A009",x"4429",x"A00A",x"4420",x"A00A",x"428E",x"A00B",x"9FD7",x"4444",x"A00A",x"A00F",x"9001",x"A000",x"4429",x"A00A",x"4420", -- 05D0-05DF 
  x"A00A",x"4280",x"440B",x"A003",x"FF83",x"32E1",x"0004",x"4784",x"42D9",x"2F0C",x"A00A",x"2F0B",x"A009",x"2F0C",x"A00A",x"426D", -- 05E0-05EF 
  x"42F0",x"4287",x"2F0C",x"A00A",x"2F0D",x"A00A",x"428E",x"A008",x"9004",x"0001",x"2F0C",x"42BB",x"8FF0",x"2F0C",x"A00A",x"2F0B", -- 05F0-05FF 
  x"A009",x"2F0C",x"A00A",x"426D",x"003C",x"4287",x"9004",x"2F0C",x"A00A",x"2F0D",x"A009",x"2F0C",x"A00A",x"426D",x"42F0",x"4287", -- 0600-060F 
  x"A00B",x"2F0C",x"A00A",x"2F0D",x"A00A",x"428E",x"A008",x"9004",x"0001",x"2F0C",x"42BB",x"8FE5",x"2F0B",x"A00A",x"2F0C",x"A00A", -- 0610-061F 
  x"B502",x"4280",x"B501",x"9003",x"0001",x"2F0C",x"42BB",x"42C6",x"B300",x"A003",x"FFBA",x"32E6",x"0002",x"4784",x"42D9",x"B502", -- 0620-062F 
  x"42F0",x"4280",x"9007",x"42C6",x"B300",x"B300",x"B300",x"B300",x"0000",x"8023",x"42C6",x"B300",x"B412",x"0000",x"B603",x"4280", -- 0630-063F 
  x"9016",x"42D9",x"42D9",x"B502",x"426D",x"B502",x"426D",x"4280",x"9004",x"B300",x"B300",x"0000",x"0000",x"B501",x"9004",x"4279", -- 0640-064F 
  x"B412",x"4279",x"B412",x"42C6",x"42C6",x"4279",x"8FE7",x"B200",x"B300",x"9002",x"FFFF",x"8001",x"0000",x"A003",x"FFCC",x"32E9", -- 0650-065F 
  x"0004",x"4784",x"42D9",x"42D9",x"0000",x"2F11",x"A00A",x"2F01",x"A00A",x"9003",x"B501",x"A00A",x"A007",x"B501",x"4279",x"B501", -- 0660-066F 
  x"A00A",x"B412",x"4279",x"A00A",x"42C6",x"42C6",x"B603",x"42D9",x"42D9",x"462E",x"9003",x"B412",x"A00D",x"B412",x"B502",x"A00D", -- 0670-067F 
  x"B502",x"A00A",x"A00D",x"A00B",x"A008",x"B502",x"B501",x"A00A",x"A007",x"2F11",x"A00A",x"4287",x"A00B",x"A008",x"9004",x"B501", -- 0680-068F 
  x"A00A",x"A007",x"8FDA",x"42C6",x"B300",x"42C6",x"B434",x"A00D",x"9004",x"B300",x"B300",x"0000",x"0000",x"A003",x"FFC0",x"32EE", -- 0690-069F 
  x"0004",x"4784",x"B412",x"0003",x"A007",x"B412",x"A003",x"FFF7",x"32F3",x"0008",x"4784",x"4047",x"4000",x"A007",x"42F9",x"A003", -- 06A0-06AF 
  x"FFF7",x"32FC",x"0006",x"4784",x"43E6",x"2F0F",x"A00A",x"2F11",x"A00A",x"B502",x"4280",x"42F9",x"2F11",x"A009",x"0020",x"45E8", -- 06B0-06BF 
  x"41B2",x"0001",x"2F01",x"A009",x"A003",x"FFEB",x"3303",x"0009",x"4784",x"2F0A",x"A00A",x"42D9",x"2F0B",x"A00A",x"42D9",x"2F0C", -- 06C0-06CF 
  x"A00A",x"42D9",x"2F0D",x"A00A",x"42D9",x"B502",x"A007",x"2F0D",x"A009",x"B501",x"2F0A",x"A009",x"B501",x"2F0B",x"A009",x"2F0C", -- 06D0-06DF 
  x"A009",x"0020",x"45E8",x"B501",x"901F",x"B603",x"4662",x"B501",x"9009",x"42D9",x"42D9",x"B200",x"42C6",x"42C6",x"46A2",x"B300", -- 06E0-06EF 
  x"4304",x"8011",x"B200",x"B603",x"456B",x"9005",x"B200",x"B300",x"0003",x"43C2",x"8008",x"B434",x"B300",x"B412",x"B300",x"2F10", -- 06F0-06FF 
  x"A00A",x"9001",x"4051",x"8FDD",x"B200",x"42C6",x"2F0D",x"A009",x"42C6",x"2F0C",x"A009",x"42C6",x"2F0B",x"A009",x"42C6",x"2F0A", -- 0700-070F 
  x"A009",x"A003",x"FFB3",x"330D",x"0004",x"4784",x"2F02",x"A00A",x"2802",x"A009",x"2F00",x"A00A",x"9006",x"003C",x"4316",x"3312", -- 0710-071F 
  x"0004",x"41EB",x"8003",x"3317",x"0002",x"41EB",x"436D",x"2F09",x"A00A",x"0100",x"44D6",x"B502",x"A00A",x"003C",x"4287",x"9002", -- 0720-072F 
  x"B200",x"802B",x"2F00",x"A00A",x"900C",x"003C",x"4316",x"331A",x"0003",x"41EB",x"46C9",x"003C",x"4316",x"331E",x"0004",x"41EB", -- 0730-073F 
  x"801C",x"001B",x"4316",x"005B",x"4316",x"0033",x"4316",x"0036",x"4316",x"006D",x"4316",x"46C9",x"2F10",x"A00A",x"A00D",x"9003", -- 0740-074F 
  x"3323",x"0002",x"41EB",x"001B",x"4316",x"005B",x"4316",x"0033",x"4316",x"0039",x"4316",x"006D",x"4316",x"8FC8",x"A003",x"FFB3", -- 0750-075F 
  x"3326",x"0005",x"4784",x"332C",x"000B",x"41EB",x"436D",x"436D",x"4716",x"A003",x"FFF5",x"3338",x"0006",x"4784",x"0000",x"2F01", -- 0760-076F 
  x"A009",x"A003",x"FFF8",x"333F",x"000C",x"4784",x"42C6",x"42D9",x"A003",x"FFF9",x"334C",x"000A",x"4784",x"42C6",x"46AB",x"A003", -- 0770-077F 
  x"FFF9",x"3357",x"0003",x"4784",x"42C6",x"2F10",x"A00A",x"9002",x"46AB",x"8001",x"42D9",x"A003",x"FFF4",x"335B",x"000A",x"4784", -- 0780-078F 
  x"46B4",x"0001",x"2F10",x"A009",x"4775",x"A003",x"FFF6",x"3366",x"0008",x"4784",x"46B4",x"0001",x"2F10",x"A009",x"477C",x"A003", -- 0790-079F 
  x"FFF6",x"336F",x"0001",x"4784",x"46B4",x"0001",x"2F10",x"A009",x"4783",x"A003",x"FFF6",x"3371",x"0001",x"4776",x"0000",x"2F10", -- 07A0-07AF 
  x"A009",x"43EF",x"4047",x"A003",x"42F9",x"476E",x"A003",x"FFF3",x"3373",x"0003",x"4784",x"2F16",x"A00A",x"9005",x"431D",x"B300", -- 07B0-07BF 
  x"431D",x"B300",x"8006",x"431D",x"4327",x"4316",x"431D",x"4327",x"4316",x"431D",x"4327",x"4316",x"431D",x"4327",x"4316",x"B300", -- 07C0-07CF 
  x"A003",x"FFE6",x"3377",x"0003",x"4784",x"337B",x"0001",x"41EB",x"0022",x"4316",x"47BB",x"0022",x"4316",x"337D",x"0001",x"41EB", -- 07D0-07DF 
  x"A003",x"FFF0",x"337F",x"0005",x"4784",x"2F16",x"A009",x"2F00",x"A00A",x"42D9",x"0000",x"2F00",x"A009",x"3385",x"0008",x"41E5", -- 07E0-07EF 
  x"46C9",x"4047",x"4000",x"A007",x"0010",x"A009",x"436D",x"003C",x"4316",x"338E",x"0006",x"41EB",x"436D",x"3395",x"0002",x"41EB", -- 07F0-07FF 
  x"0000",x"B603",x"A007",x"B501",x"2F03",x"4287",x"9002",x"B300",x"2F04",x"B501",x"2F17",x"4287",x"9005",x"B300",x"2F00",x"2F80", -- 0800-080F 
  x"A009",x"2F80",x"A00A",x"47D5",x"4279",x"B501",x"0010",x"4287",x"9FE8",x"B300",x"3398",x"0004",x"41EB",x"B501",x"4346",x"339D", -- 0810-081F 
  x"0001",x"41EB",x"B501",x"000F",x"A007",x"4360",x"0010",x"A007",x"B603",x"42A0",x"A00B",x"9FD0",x"B200",x"436D",x"003C",x"4316", -- 0820-082F 
  x"339F",x"0007",x"41EB",x"42C6",x"2F00",x"A009",x"A003",x"FFAA",x"33A7",x"0005",x"4060",x"2F20",x"FFFB",x"33AD",x"0008",x"4784", -- 0830-083F 
  x"2F20",x"A00A",x"B501",x"406B",x"B501",x"4279",x"2F20",x"A009",x"A009",x"A003",x"FFF2",x"33B6",x"0004",x"4784",x"B501",x"900D", -- 0840-084F 
  x"42D9",x"B502",x"A00A",x"B502",x"A009",x"B412",x"4279",x"B412",x"4279",x"42C6",x"0001",x"4280",x"8FF1",x"B300",x"B200",x"A003", -- 0850-085F 
  x"FFEA",x"33BB",x"0004",x"4784",x"B434",x"B434",x"B501",x"9009",x"42D9",x"B603",x"A009",x"0001",x"A007",x"42C6",x"0001",x"4280", -- 0860-086F 
  x"8FF5",x"B300",x"B200",x"A003",x"FFEC",x"33C0",x"0004",x"4784",x"B412",x"B501",x"A00A",x"4360",x"0001",x"A007",x"B412",x"0001", -- 0870-087F 
  x"4280",x"B501",x"A00D",x"9FF4",x"B300",x"A003",x"FFEE",x"33C5",x"0003",x"4784",x"B603",x"428E",x"9001",x"B412",x"B300",x"A003", -- 0880-088F 
  x"FFF6",x"33C9",x"0003",x"4784",x"B603",x"42A0",x"9001",x"B412",x"B300",x"A003",x"FFF6",x"33CD",x"0003",x"4784",x"B501",x"A00F", -- 0890-089F 
  x"9001",x"A000",x"A003",x"FFF7",x"33D1",x"0006",x"410A",x"A017",x"A003",x"FFFA",x"33D8",x"0007",x"410A",x"A018",x"A003",x"FFFA", -- 08A0-08AF 
  x"33E0",x"0009",x"4784",x"42D9",x"A017",x"A018",x"9FFD",x"42C6",x"B300",x"A003",x"FFF5",x"33EA",x"0001",x"4060",x"1401",x"FFFB", -- 08B0-08BF 
  x"33EC",x"0001",x"4060",x"1601",x"FFFB",x"33EE",x"0001",x"4060",x"1801",x"FFFB",x"33F0",x"0004",x"4784",x"0007",x"43FC",x"444D", -- 08C0-08CF 
  x"A009",x"4444",x"A009",x"443B",x"A009",x"4432",x"A009",x"4429",x"A009",x"4420",x"A009",x"4417",x"A009",x"4417",x"A00A",x"4432", -- 08D0-08DF 
  x"A00A",x"9001",x"A00B",x"4420",x"A00A",x"443B",x"A00A",x"A007",x"4279",x"444D",x"A00A",x"B502",x"0000",x"4864",x"444D",x"A00A", -- 08E0-08EF 
  x"B501",x"4429",x"A00A",x"4420",x"A00A",x"0000",x"B60C",x"A00A",x"B434",x"B434",x"4444",x"A00A",x"443B",x"A00A",x"48B3",x"B300", -- 08F0-08FF 
  x"A009",x"B300",x"B434",x"0001",x"A007",x"B434",x"0001",x"A007",x"B434",x"FFFF",x"A007",x"B501",x"A00D",x"9FE7",x"B300",x"B200", -- 0900-090F 
  x"440B",x"A003",x"FFB7",x"33F5",x"0006",x"4784",x"0007",x"43FC",x"444D",x"A009",x"4444",x"A009",x"443B",x"A009",x"4432",x"A009", -- 0910-091F 
  x"4429",x"A009",x"4420",x"A009",x"4417",x"A009",x"4417",x"A00A",x"4420",x"A00A",x"443B",x"A00A",x"488A",x"4279",x"444D",x"A00A", -- 0920-092F 
  x"4417",x"A00A",x"4432",x"A00A",x"4287",x"903C",x"0000",x"4420",x"A00A",x"443B",x"A00A",x"488A",x"0000",x"B434",x"B502",x"B501", -- 0930-093F 
  x"4420",x"A00A",x"428E",x"9009",x"4429",x"A00A",x"B501",x"A00A",x"B412",x"4279",x"4429",x"A009",x"8001",x"0000",x"B412",x"443B", -- 0940-094F 
  x"A00A",x"428E",x"9009",x"4444",x"A00A",x"B501",x"A00A",x"B412",x"4279",x"4444",x"A009",x"8001",x"0000",x"A001",x"444D",x"A00A", -- 0950-095F 
  x"B501",x"4279",x"444D",x"A009",x"A009",x"B434",x"B434",x"0001",x"A007",x"B603",x"4280",x"A00D",x"9FD0",x"B200",x"444D",x"A00A", -- 0960-096F 
  x"A009",x"8065",x"B412",x"0001",x"4280",x"B412",x"0001",x"4420",x"A00A",x"443B",x"A00A",x"488A",x"0000",x"B434",x"B502",x"B501", -- 0970-097F 
  x"4420",x"A00A",x"428E",x"9009",x"4429",x"A00A",x"B501",x"A00A",x"B412",x"4279",x"4429",x"A009",x"8001",x"0000",x"B412",x"443B", -- 0980-098F 
  x"A00A",x"428E",x"900A",x"4444",x"A00A",x"B501",x"A00A",x"B412",x"4279",x"4444",x"A009",x"A00B",x"8001",x"FFFF",x"A001",x"444D", -- 0990-099F 
  x"A00A",x"B501",x"4279",x"444D",x"A009",x"A009",x"B434",x"B434",x"0001",x"A007",x"B603",x"4280",x"A00D",x"9FCF",x"B200",x"A00D", -- 09A0-09AF 
  x"9026",x"B501",x"444D",x"A009",x"B434",x"A00B",x"B434",x"B434",x"0001",x"4420",x"A00A",x"443B",x"A00A",x"488A",x"0000",x"B434", -- 09B0-09BF 
  x"0000",x"444D",x"A00A",x"A00A",x"A00B",x"A001",x"444D",x"A00A",x"B501",x"4279",x"444D",x"A009",x"A009",x"B434",x"B434",x"0001", -- 09C0-09CF 
  x"A007",x"B603",x"4280",x"A00D",x"9FEA",x"B200",x"B300",x"440B",x"A003",x"FF39",x"33FC",x"0004",x"410A",x"A014",x"A003",x"FFFA", -- 09D0-09DF 
  x"3401",x"0005",x"4784",x"0010",x"42D9",x"A014",x"42C6",x"0001",x"4280",x"B501",x"A00D",x"9FF8",x"B200",x"A003",x"FFF1",x"3407", -- 09E0-09EF 
  x"0004",x"4784",x"0000",x"B434",x"B434",x"49E3",x"A003",x"FFF7",x"340C",x"0004",x"4784",x"B502",x"A00F",x"9012",x"B412",x"A000", -- 09F0-09FF 
  x"B412",x"B501",x"A00F",x"9006",x"A000",x"49F2",x"B412",x"A000",x"B412",x"8005",x"49F2",x"A000",x"B412",x"A000",x"B412",x"8008", -- 0A00-0A0F 
  x"B501",x"A00F",x"9004",x"A000",x"49F2",x"A000",x"8001",x"49F2",x"A003",x"FFDE",x"3411",x"0001",x"4784",x"49FB",x"B412",x"B300", -- 0A10-0A1F 
  x"A003",x"FFF8",x"3413",x"0003",x"4784",x"49FB",x"B300",x"A003",x"FFF9",x"3417",x"0004",x"4784",x"0007",x"43FC",x"444D",x"A009", -- 0A20-0A2F 
  x"4444",x"A009",x"443B",x"A009",x"4432",x"A009",x"4429",x"A009",x"4420",x"A009",x"4417",x"A009",x"4420",x"A00A",x"443B",x"A00A", -- 0A30-0A3F 
  x"428E",x"900A",x"4417",x"A00A",x"4420",x"A00A",x"4429",x"A00A",x"0000",x"0000",x"0000",x"80E1",x"4420",x"A00A",x"0000",x"4429", -- 0A40-0A4F 
  x"A00A",x"B502",x"A007",x"A00A",x"A00B",x"B502",x"444D",x"A00A",x"A007",x"A009",x"0001",x"A007",x"B603",x"4280",x"A00D",x"9FEF", -- 0A50-0A5F 
  x"B200",x"444D",x"A00A",x"4420",x"A00A",x"A007",x"443B",x"A00A",x"4280",x"4429",x"A009",x"FFFF",x"444D",x"A00A",x"4420",x"A00A", -- 0A60-0A6F 
  x"A007",x"A009",x"0001",x"4420",x"42BB",x"4420",x"A00A",x"443B",x"A00A",x"4280",x"0000",x"4429",x"A00A",x"443B",x"A00A",x"A007", -- 0A70-0A7F 
  x"A00A",x"A00B",x"4429",x"A00A",x"443B",x"A00A",x"A007",x"0001",x"4280",x"A00A",x"A00B",x"4444",x"A00A",x"443B",x"A00A",x"A007", -- 0A80-0A8F 
  x"0001",x"4280",x"A00A",x"49E3",x"B412",x"B300",x"B501",x"4429",x"A00A",x"443B",x"A00A",x"A007",x"4279",x"A009",x"0000",x"4429", -- 0A90-0A9F 
  x"A00A",x"4444",x"A00A",x"443B",x"A00A",x"48B3",x"B200",x"B412",x"B300",x"0000",x"4429",x"A00A",x"443B",x"A00A",x"A007",x"A00A", -- 0AA0-0AAF 
  x"A001",x"4429",x"A00A",x"443B",x"A00A",x"A007",x"A009",x"902C",x"0001",x"443B",x"A00A",x"0000",x"B434",x"B502",x"4429",x"A00A", -- 0AB0-0ABF 
  x"B502",x"A007",x"A00A",x"B412",x"4444",x"A00A",x"A007",x"A00A",x"A00B",x"A001",x"B412",x"42D9",x"B502",x"4429",x"A00A",x"A007", -- 0AC0-0ACF 
  x"A009",x"42C6",x"B434",x"B434",x"0001",x"A007",x"B603",x"4280",x"A00D",x"9FE2",x"B200",x"FFFF",x"4429",x"A00A",x"443B",x"A00A", -- 0AD0-0ADF 
  x"A007",x"4279",x"42BB",x"8FD3",x"FFFF",x"4429",x"42BB",x"0001",x"A007",x"B603",x"4280",x"A00D",x"9F8E",x"B200",x"443B",x"A00A", -- 0AE0-0AEF 
  x"0000",x"444D",x"A00A",x"B502",x"A007",x"A00A",x"A00B",x"B502",x"444D",x"A00A",x"A007",x"A009",x"0001",x"A007",x"B603",x"4280", -- 0AF0-0AFF 
  x"A00D",x"9FEF",x"B200",x"443B",x"A00A",x"444D",x"A00A",x"0001",x"4280",x"A009",x"4420",x"A00A",x"443B",x"A00A",x"4280",x"444D", -- 0B00-0B0F 
  x"A00A",x"443B",x"A00A",x"A007",x"A009",x"4417",x"A00A",x"443B",x"A00A",x"444D",x"A00A",x"4417",x"A00A",x"4432",x"A00A",x"9001", -- 0B10-0B1F 
  x"A00B",x"4420",x"A00A",x"443B",x"A00A",x"4280",x"444D",x"A00A",x"443B",x"A00A",x"A007",x"0001",x"A007",x"440B",x"A003",x"FEF9", -- 0B20-0B2F 
  x"341C",x"0008",x"4060",x"2F21",x"FFFB",x"3425",x"0008",x"4060",x"2F22",x"FFFB",x"342E",x"0008",x"4060",x"2F23",x"FFFB",x"3437", -- 0B30-0B3F 
  x"000E",x"4060",x"2F24",x"FFFB",x"3446",x"000C",x"4060",x"2F25",x"FFFB",x"3453",x"0006",x"4060",x"2F26",x"FFFB",x"345A",x"000D", -- 0B40-0B4F 
  x"4784",x"B502",x"A00D",x"9004",x"B200",x"B300",x"0000",x"8031",x"B603",x"A007",x"0001",x"4280",x"B501",x"A00A",x"A00D",x"A00B", -- 0B50-0B5F 
  x"9FF9",x"0001",x"A007",x"B502",x"488A",x"B603",x"4287",x"9004",x"B200",x"B200",x"0000",x"801D",x"B502",x"4280",x"B502",x"A00A", -- 0B60-0B6F 
  x"C000",x"A008",x"A00D",x"B502",x"0001",x"4287",x"A008",x"9003",x"B300",x"A00A",x"8009",x"B502",x"0001",x"4280",x"A009",x"0001", -- 0B70-0B7F 
  x"4280",x"4047",x"4000",x"A00E",x"B412",x"B300",x"B412",x"9001",x"A000",x"A003",x"FFC3",x"3468",x"000C",x"4784",x"B501",x"A00A", -- 0B80-0B8F 
  x"B501",x"A00F",x"9003",x"A000",x"FFFF",x"8001",x"0000",x"B434",x"B434",x"B501",x"4047",x"4000",x"A008",x"9009",x"B412",x"B300", -- 0B90-0B9F 
  x"3FFF",x"A008",x"B501",x"A00A",x"B412",x"4279",x"8004",x"B502",x"A009",x"0001",x"B412",x"A003",x"FFDE",x"3475",x"000B",x"4784", -- 0BA0-0BAF 
  x"2F23",x"A00A",x"B603",x"A009",x"4279",x"B603",x"A007",x"2F23",x"A009",x"B603",x"B412",x"0000",x"4864",x"B412",x"B300",x"2F23", -- 0BB0-0BBF 
  x"A00A",x"2F25",x"A00A",x"428E",x"A00B",x"9002",x"0369",x"43C2",x"A003",x"FFE3",x"3481",x"0010",x"4784",x"2F22",x"A009",x"2F21", -- 0BC0-0BCF 
  x"A009",x"2F21",x"4B8E",x"B502",x"42D9",x"2F22",x"4B8E",x"B502",x"42C6",x"A007",x"4279",x"4BB0",x"A003",x"FFEC",x"3492",x"0002", -- 0BD0-0BDF 
  x"4784",x"4BCD",x"4916",x"4B51",x"A003",x"FFF8",x"3495",x"0002",x"4784",x"A000",x"4BE1",x"A003",x"FFF9",x"3498",x"0002",x"4784", -- 0BE0-0BEF 
  x"4BCD",x"48CD",x"4B51",x"A003",x"FFF8",x"349B",x"0007",x"4776",x"2F11",x"A00A",x"0004",x"A007",x"46AB",x"A003",x"FFF6",x"34A3", -- 0BF0-0BFF 
  x"0005",x"4784",x"B501",x"A00D",x"9002",x"0000",x"43C2",x"B501",x"2F21",x"A009",x"2F21",x"4B8E",x"B434",x"B300",x"B502",x"A007", -- 0C00-0C0F 
  x"0001",x"4280",x"A00A",x"B412",x"0001",x"42A0",x"9018",x"0001",x"B502",x"A00F",x"A00B",x"9007",x"B412",x"B501",x"A007",x"B412", -- 0C10-0C1F 
  x"B501",x"4BE1",x"8FF5",x"B412",x"B300",x"B501",x"2F26",x"A009",x"B434",x"B502",x"4BF0",x"B434",x"B434",x"4BF0",x"8004",x"B300", -- 0C20-0C2F 
  x"0001",x"2F26",x"A009",x"4BCD",x"4A2C",x"4B51",x"42D9",x"4B51",x"42C6",x"2F26",x"A00A",x"0001",x"4280",x"9007",x"B412",x"2F26", -- 0C30-0C3F 
  x"A00A",x"4C02",x"B412",x"B300",x"B412",x"A003",x"FFB8",x"34A9",x"0004",x"4784",x"0000",x"42D9",x"431D",x"B501",x"9007",x"4327", -- 0C40-0C4F 
  x"4316",x"42C6",x"B300",x"FFFF",x"42D9",x"8001",x"B300",x"431D",x"B501",x"42F0",x"A00E",x"9007",x"4327",x"4316",x"42C6",x"B300", -- 0C50-0C5F 
  x"FFFF",x"42D9",x"8001",x"B300",x"431D",x"B501",x"42F0",x"A00E",x"9003",x"4327",x"4316",x"8001",x"B300",x"431D",x"4327",x"4316", -- 0C60-0C6F 
  x"B300",x"42C6",x"B300",x"A003",x"FFD2",x"34AE",x"0002",x"4784",x"2F21",x"A009",x"2F21",x"4B8E",x"B434",x"9003",x"34B1",x"0001", -- 0C70-0C7F 
  x"41EB",x"B502",x"A007",x"0001",x"4280",x"B501",x"A00A",x"4C4A",x"B412",x"0001",x"4280",x"B412",x"B502",x"900A",x"0001",x"4280", -- 0C80-0C8F 
  x"B501",x"A00A",x"4346",x"B412",x"0001",x"4280",x"B412",x"8FF4",x"B300",x"B300",x"0020",x"4316",x"A003",x"FFD7",x"34B3",x"0003", -- 0C90-0C9F 
  x"4784",x"B412",x"4C78",x"4C78",x"A003",x"FFF8",x"34B7",x"000B",x"4060",x"2F27",x"FFFB",x"34C3",x"0009",x"4060",x"2F28",x"FFFB", -- 0CA0-0CAF 
  x"34CD",x"000D",x"4784",x"2F23",x"A00A",x"A003",x"FFF9",x"34DB",x"000D",x"4784",x"2F23",x"A009",x"A003",x"FFF9",x"34E9",x"000B", -- 0CB0-0CBF 
  x"4784",x"2F28",x"A00A",x"2F27",x"A009",x"2F23",x"A00A",x"2F28",x"A009",x"A003",x"FFF3",x"34F5",x"0004",x"4784",x"2F24",x"A00A", -- 0CC0-0CCF 
  x"2F23",x"A009",x"4CC1",x"4CC1",x"A003",x"FFF5",x"34FA",x"0003",x"4784",x"B501",x"2F21",x"A009",x"2F21",x"4B8E",x"B501",x"2F21", -- 0CD0-0CDF 
  x"4280",x"B300",x"0001",x"901A",x"B502",x"2F23",x"A00A",x"4279",x"B412",x"484E",x"2F23",x"A00A",x"4279",x"B502",x"4279",x"2F23", -- 0CE0-0CEF 
  x"42BB",x"2F23",x"A00A",x"2F25",x"A00A",x"428E",x"A00B",x"9002",x"0369",x"43C2",x"4B51",x"B412",x"B300",x"8002",x"B200",x"B300", -- 0CF0-0CFF 
  x"A003",x"FFD4",x"34FE",x"0003",x"4784",x"B412",x"4CD9",x"B412",x"4CD9",x"A003",x"FFF7",x"3502",x"0002",x"4784",x"4CB3",x"B434", -- 0D00-0D0F 
  x"B434",x"4C02",x"B412",x"B300",x"B412",x"4CBA",x"4CD9",x"A003",x"FFF2",x"3505",x"0004",x"4784",x"4CB3",x"B434",x"B434",x"4C02", -- 0D10-0D1F 
  x"B300",x"B412",x"4CBA",x"4CD9",x"A003",x"FFF3",x"350A",x"0004",x"4784",x"4CB3",x"B434",x"B434",x"B501",x"9004",x"B412",x"B502", -- 0D20-0D2F 
  x"4D1C",x"8FFA",x"B300",x"B412",x"4CBA",x"4CD9",x"A003",x"FFEE",x"350F",x"0003",x"4784",x"4CB3",x"B434",x"B434",x"B603",x"4D29", -- 0D30-0D3F 
  x"B434",x"B502",x"4D0E",x"B434",x"B434",x"4D0E",x"B434",x"4CBA",x"4D05",x"A003",x"FFED",x"3513",x"0007",x"4784",x"4CB3",x"B434", -- 0D40-0D4F 
  x"B434",x"0007",x"43FC",x"4420",x"A009",x"4417",x"A009",x"0000",x"4420",x"A00A",x"9063",x"B501",x"4429",x"A009",x"0001",x"4444", -- 0D50-0D5F 
  x"A009",x"FFFF",x"444D",x"A009",x"4417",x"A00A",x"4429",x"A00A",x"A007",x"426D",x"002B",x"4287",x"9009",x"4429",x"A00A",x"4279", -- 0D60-0D6F 
  x"4429",x"A009",x"0000",x"444D",x"A009",x"8016",x"4417",x"A00A",x"4429",x"A00A",x"A007",x"426D",x"002D",x"4287",x"900D",x"4429", -- 0D70-0D7F 
  x"A00A",x"4279",x"4429",x"A009",x"0000",x"444D",x"A009",x"4444",x"A00A",x"A000",x"4444",x"A009",x"444D",x"A00A",x"9FD2",x"4429", -- 0D80-0D8F 
  x"A00A",x"4420",x"A00A",x"428E",x"9029",x"4417",x"A00A",x"4429",x"A00A",x"A007",x"426D",x"B501",x"9015",x"4542",x"A00B",x"9007", -- 0D90-0D9F 
  x"B300",x"4420",x"A00A",x"A000",x"4420",x"A009",x"800A",x"B412",x"2F08",x"A00A",x"4BF0",x"4BE1",x"4429",x"A00A",x"4279",x"4429", -- 0DA0-0DAF 
  x"A009",x"8005",x"B300",x"4429",x"A00A",x"4420",x"A009",x"4429",x"A00A",x"4420",x"A00A",x"428E",x"A00B",x"9FD7",x"4444",x"A00A", -- 0DB0-0DBF 
  x"A00F",x"9001",x"A000",x"4429",x"A00A",x"4420",x"A00A",x"4280",x"B501",x"9006",x"B300",x"4417",x"A00A",x"4429",x"A00A",x"A007", -- 0DC0-0DCF 
  x"440B",x"B434",x"4CBA",x"B412",x"4CD9",x"B412",x"A003",x"FF73",x"351B",x"0002",x"0022",x"41CA",x"4D4E",x"B300",x"A003",x"FFF8", -- 0DD0-0DDF 
  x"351E",x"0002",x"4784",x"4CB3",x"B434",x"B434",x"0004",x"43FC",x"B501",x"A00F",x"9002",x"0012",x"43C2",x"0002",x"4432",x"A009", -- 0DE0-0DEF 
  x"4429",x"A009",x"4420",x"A009",x"0001",x"4429",x"A00A",x"4432",x"A00A",x"49FB",x"4429",x"A009",x"9003",x"4420",x"A00A",x"4BF0", -- 0DF0-0DFF 
  x"4429",x"A00A",x"9008",x"4420",x"A00A",x"4420",x"A00A",x"4BF0",x"4420",x"A009",x"8FEA",x"440B",x"B412",x"4CBA",x"4CD9",x"A003", -- 0E00-0E0F 
  x"FFCF",x"3521",x"0002",x"4784",x"2F08",x"A00A",x"0010",x"4287",x"9002",x"4C78",x"802C",x"4CB3",x"B412",x"B501",x"A00F",x"9004", -- 0E10-0E1F 
  x"A000",x"3524",x"0001",x"41EB",x"B501",x"A00D",x"9005",x"3526",x"0002",x"41EB",x"B300",x"801A",x"FFFF",x"B412",x"B501",x"9004", -- 0E20-0E2F 
  x"2F08",x"A00A",x"4C02",x"8FFA",x"B300",x"B501",x"A00F",x"A00B",x"900A",x"0030",x"A007",x"B501",x"0039",x"42A0",x"9002",x"0007", -- 0E30-0E3F 
  x"A007",x"4316",x"8FF2",x"0020",x"4316",x"B300",x"4CBA",x"A003",x"FFC8",x"3529",x"0003",x"4784",x"B412",x"4E14",x"4E14",x"A003", -- 0E40-0E4F 
  x"FFF8",x"352D",x"0006",x"4784",x"3FFF",x"A008",x"B501",x"4279",x"B412",x"A00A",x"A003",x"FFF5",x"3534",x"0004",x"4784",x"489E", -- 0E50-0E5F 
  x"B501",x"4047",x"4000",x"428E",x"9003",x"B300",x"0000",x"800A",x"4E54",x"B412",x"B300",x"4047",x"4000",x"428E",x"9002",x"0000", -- 0E60-0E6F 
  x"8001",x"FFFF",x"A003",x"FFE8",x"3539",x"0001",x"4784",x"B502",x"4E5F",x"9011",x"B412",x"4E54",x"3FFF",x"A008",x"B434",x"B603", -- 0E70-0E7F 
  x"42A0",x"9005",x"B412",x"B300",x"A007",x"A00A",x"8003",x"B200",x"B300",x"0000",x"8003",x"9002",x"B300",x"0000",x"A003",x"FFE4", -- 0E80-0E8F 
  x"353B",x"0001",x"4784",x"B603",x"4E77",x"A003",x"FFF9",x"353D",x"0001",x"4784",x"B501",x"42D9",x"B434",x"B434",x"B502",x"4E5F", -- 0E90-0E9F 
  x"A00D",x"B502",x"A00D",x"A008",x"42C6",x"4E5F",x"A00D",x"A008",x"9002",x"B200",x"806F",x"B502",x"4E5F",x"A00D",x"9017",x"B501", -- 0EA0-0EAF 
  x"4279",x"4BB0",x"B434",x"B502",x"A009",x"4047",x"4000",x"B502",x"0001",x"4280",x"42BB",x"B501",x"42D9",x"A007",x"A009",x"42C6", -- 0EB0-0EBF 
  x"0001",x"4280",x"4047",x"4000",x"A007",x"8054",x"B502",x"4E54",x"3FFF",x"A008",x"B434",x"B603",x"42A0",x"9008",x"B412",x"B300", -- 0EC0-0ECF 
  x"B434",x"42D9",x"A007",x"A009",x"42C6",x"801B",x"B501",x"4279",x"4BB0",x"B412",x"42D9",x"B501",x"42D9",x"B412",x"484E",x"B300", -- 0ED0-0EDF 
  x"42C6",x"4047",x"4000",x"B502",x"0001",x"4280",x"42BB",x"B412",x"B502",x"42C6",x"A007",x"A009",x"0001",x"4280",x"4047",x"4000", -- 0EE0-0EEF 
  x"A007",x"4E54",x"3FFF",x"A008",x"B603",x"A007",x"0001",x"4280",x"A00A",x"A00D",x"B502",x"0001",x"42A0",x"A008",x"9003",x"0001", -- 0EF0-0EFF 
  x"4280",x"8FF2",x"B502",x"A00A",x"4E5F",x"A00D",x"B502",x"0001",x"4287",x"A008",x"9003",x"B300",x"A00A",x"800C",x"B412",x"0001", -- 0F00-0F0F 
  x"4280",x"B412",x"4047",x"4000",x"A007",x"B502",x"A009",x"4047",x"4000",x"A007",x"A003",x"FF7B",x"353F",x"0002",x"4784",x"B501", -- 0F10-0F1F 
  x"4E5F",x"9017",x"3542",x"0002",x"41EB",x"4E54",x"3FFF",x"A008",x"B502",x"A007",x"B412",x"B603",x"42A0",x"9006",x"B501",x"A00A", -- 0F20-0F2F 
  x"4F1F",x"0001",x"A007",x"8FF7",x"B200",x"3545",x"0002",x"41EB",x"8001",x"4E14",x"A003",x"FFE0",x"3548",x"0006",x"4060",x"2F29", -- 0F30-0F3F 
  x"FFFB",x"354F",x"0001",x"4784",x"2F29",x"A00A",x"2801",x"A00A",x"2F29",x"A009",x"A003",x"FFF5",x"3551",x"0001",x"4784",x"0000", -- 0F40-0F4F 
  x"2801",x"A00A",x"0001",x"4280",x"2F29",x"A00A",x"4280",x"900A",x"2801",x"A00A",x"0002",x"4280",x"2F29",x"A00A",x"4280",x"B434", -- 0F50-0F5F 
  x"4E9A",x"8FEE",x"B412",x"2F29",x"A009",x"A003",x"FFE5",x"3553",x"0005",x"4784",x"B501",x"4E5F",x"901C",x"B501",x"42D9",x"4E54", -- 0F60-0F6F 
  x"3FFF",x"A008",x"B412",x"B502",x"A007",x"FFFF",x"A007",x"B412",x"B501",x"900C",x"B412",x"B501",x"A00A",x"4F6A",x"B502",x"A009", -- 0F70-0F7F 
  x"FFFF",x"A007",x"B412",x"FFFF",x"A007",x"8FF2",x"B200",x"42C6",x"8001",x"4CD9",x"A003",x"FFDB",x"3559",x"0007",x"4784",x"B501", -- 0F80-0F8F 
  x"4E5F",x"902A",x"4E54",x"3FFF",x"A008",x"B501",x"9023",x"B412",x"436D",x"B502",x"4360",x"B501",x"4360",x"B501",x"A00A",x"B501", -- 0F90-0F9F 
  x"4360",x"B501",x"489E",x"4047",x"4000",x"428E",x"9005",x"FFFF",x"4360",x"FFFF",x"4360",x"8005",x"B501",x"489E",x"4E54",x"4360", -- 0FA0-0FAF 
  x"4360",x"B501",x"4F1F",x"4F8F",x"0001",x"A007",x"B412",x"FFFF",x"A007",x"8FDB",x"B200",x"8001",x"B300",x"A003",x"FFCD",x"3561", -- 0FB0-0FBF 
  x"000B",x"4784",x"0008",x"43FC",x"4CB3",x"4417",x"A009",x"4420",x"A009",x"0001",x"4420",x"A00A",x"4429",x"A009",x"FFFF",x"4429", -- 0FC0-0FCF 
  x"42BB",x"4456",x"A009",x"0000",x"4444",x"A009",x"0000",x"444D",x"A009",x"B501",x"4429",x"A00A",x"4E77",x"4429",x"A00A",x"4E77", -- 0FD0-0FDF 
  x"4420",x"A00A",x"4432",x"A009",x"FFFF",x"4432",x"42BB",x"B502",x"4432",x"A00A",x"4E77",x"4429",x"A00A",x"4E77",x"4444",x"A00A", -- 0FE0-0FEF 
  x"4432",x"A00A",x"B434",x"4E9A",x"4444",x"A009",x"B502",x"4429",x"A00A",x"4E77",x"4432",x"A00A",x"4E77",x"444D",x"A00A",x"4432", -- 0FF0-0FFF 
  x"A00A",x"B434",x"4E9A",x"444D",x"A009",x"4432",x"A00A",x"A00D",x"9FDB",x"4444",x"A00A",x"4429",x"A00A",x"4E77",x"4456",x"A00A", -- 1000-100F 
  x"4BE1",x"4444",x"A00A",x"4429",x"A00A",x"B434",x"4E9A",x"4444",x"A009",x"444D",x"A00A",x"4429",x"A00A",x"4E77",x"4456",x"A00A", -- 1010-101F 
  x"4BE9",x"444D",x"A00A",x"4429",x"A00A",x"B434",x"4E9A",x"444D",x"A009",x"4420",x"A00A",x"4432",x"A009",x"FFFF",x"4432",x"42BB", -- 1020-102F 
  x"B502",x"4432",x"A00A",x"4E77",x"4420",x"A00A",x"443B",x"A009",x"FFFF",x"443B",x"42BB",x"4CB3",x"B434",x"B434",x"B412",x"B502", -- 1030-103F 
  x"443B",x"A00A",x"4E77",x"B502",x"4BF0",x"4444",x"A00A",x"4432",x"A00A",x"4E77",x"444D",x"A00A",x"443B",x"A00A",x"4E77",x"4BF0", -- 1040-104F 
  x"4BE9",x"4456",x"A00A",x"4D0E",x"B43C",x"B412",x"4CBA",x"B412",x"4CD9",x"B412",x"443B",x"A00A",x"B434",x"4E9A",x"443B",x"A00A", -- 1050-105F 
  x"A00D",x"9FD6",x"B434",x"4432",x"A00A",x"B434",x"4E9A",x"B412",x"4432",x"A00A",x"A00D",x"9FC1",x"4CD9",x"4417",x"A00A",x"4CBA", -- 1060-106F 
  x"B412",x"4F6A",x"B412",x"4CD9",x"4429",x"A00A",x"A00D",x"9F56",x"440B",x"A003",x"FF44",x"356D",x"0011",x"4784",x"0003",x"43FC", -- 1070-107F 
  x"4417",x"A009",x"0000",x"4417",x"A00A",x"4420",x"A009",x"4420",x"A00A",x"B501",x"9023",x"0001",x"4280",x"4420",x"A009",x"4420", -- 1080-108F 
  x"A00A",x"4E93",x"4417",x"A00A",x"4429",x"A009",x"4429",x"A00A",x"B501",x"9011",x"0001",x"4280",x"4429",x"A009",x"4429",x"A00A", -- 1090-109F 
  x"4420",x"A00A",x"0001",x"A007",x"4429",x"A00A",x"0001",x"A007",x"4DE3",x"4E9A",x"8FEB",x"B300",x"4E9A",x"8FD9",x"B300",x"440B", -- 10A0-10AF 
  x"A003",x"FFC9",x"357F",x"0005",x"4784",x"2F11",x"A00A",x"B501",x"4279",x"A00A",x"B502",x"0002",x"A007",x"A00A",x"4335",x"0020", -- 10B0-10BF 
  x"4316",x"B501",x"A00A",x"9004",x"B501",x"A00A",x"A007",x"8FEF",x"B300",x"A003",x"FFE7",x"3585",x"0005",x"4784",x"2F11",x"A00A", -- 10C0-10CF 
  x"B501",x"4360",x"B501",x"4279",x"A00A",x"B502",x"0002",x"A007",x"A00A",x"4335",x"0020",x"4316",x"B501",x"A00A",x"9004",x"B501", -- 10D0-10DF 
  x"A00A",x"A007",x"8FED",x"B300",x"A003",x"FFE5",x"358B",x"0006",x"4060",x"A003",x"FFFB",x"3592",x"0008",x"4784",x"43E6",x"0020", -- 10E0-10EF 
  x"45E8",x"4662",x"B501",x"9012",x"46A2",x"B300",x"4279",x"41F1",x"B412",x"2F0F",x"A009",x"B501",x"46AB",x"4047",x"A003",x"42F9", -- 10F0-10FF 
  x"2F0F",x"A009",x"0001",x"2F10",x"A009",x"8003",x"B200",x"0003",x"43C2",x"A003",x"FFE0",x"359B",x"0006",x"4784",x"0020",x"45E8", -- 1100-110F 
  x"4662",x"900E",x"2F0F",x"A009",x"41F1",x"B501",x"A00A",x"A007",x"2F11",x"A009",x"41F1",x"4279",x"A00A",x"2F13",x"A009",x"8004", -- 1110-111F 
  x"B300",x"35A2",x"000F",x"41EB",x"A003",x"FFE5",x"35B2",x"000A",x"4784",x"436D",x"B501",x"0000",x"4287",x"9003",x"35BD",x"0013", -- 1120-112F 
  x"41EB",x"B501",x"0003",x"4287",x"9003",x"35D1",x"0014",x"41EB",x"B501",x"0006",x"4287",x"9003",x"35E6",x"0014",x"41EB",x"B501", -- 1130-113F 
  x"0009",x"4287",x"9003",x"35FB",x"0030",x"41EB",x"B501",x"0012",x"4287",x"9003",x"362C",x"0012",x"41EB",x"B501",x"0369",x"4287", -- 1140-114F 
  x"9003",x"363F",x"0013",x"41EB",x"B501",x"1234",x"4287",x"9003",x"3653",x"004C",x"41EB",x"A003",x"FFC9",x"36A0",x"0005",x"4784", -- 1150-115F 
  x"47A4",x"41F1",x"0003",x"4280",x"B501",x"4360",x"A00A",x"4279",x"B501",x"4360",x"A00A",x"B501",x"4360",x"0040",x"4280",x"41F1", -- 1160-116F 
  x"B412",x"0007",x"A008",x"2F18",x"A007",x"A009",x"A003",x"FFE5",x"36A6",x"0002",x"4784",x"0007",x"4316",x"36A9",x"0008",x"41EB", -- 1170-117F 
  x"A003",x"FFF6",x"36B2",x"0002",x"4784",x"0007",x"4316",x"36B5",x"0004",x"41EB",x"4716",x"A003",x"FFF5",x"36BA",x"0002",x"4784", -- 1180-118F 
  x"36BD",x"0029",x"41EB",x"436D",x"FA00",x"0100",x"44D6",x"46C9",x"36E7",x"0002",x"41EB",x"A003",x"FFF0",x"36EA",x"0005",x"4784", -- 1190-119F 
  x"2F09",x"A00A",x"0100",x"44D6",x"A003",x"FFF7",x"36F0",x"0007",x"4776",x"003C",x"4316",x"36F8",x"0004",x"41EB",x"436D",x"51A0", -- 11A0-11AF 
  x"36FD",x"0007",x"41E5",x"462E",x"9FF9",x"003C",x"4316",x"3705",x"0003",x"41EB",x"A003",x"FFEA",x"3709",x"0003",x"4784",x"0010", -- 11B0-11BF 
  x"2F08",x"A009",x"A003",x"FFF8",x"370D",x"0007",x"4784",x"000A",x"2F08",x"A009",x"A003",x"FFF8",x"3715",x"0005",x"4784",x"B501", -- 11C0-11CF 
  x"3FFF",x"42A0",x"B502",x"C000",x"428E",x"A00E",x"9002",x"1234",x"43C2",x"42F9",x"A003",x"51CF",x"A003",x"4D4E",x"A003",x"FFEC", -- 11D0-11DF 
  x"371B",x"0002",x"4784",x"4360",x"A003",x"FFFA",x"371E",x"0002",x"4784",x"A007",x"A003",x"FFFA",x"3721",x"0002",x"4784",x"4280", -- 11E0-11EF 
  x"A003",x"FFFA",x"3724",x"0002",x"4784",x"42A7",x"A003",x"FFFA",x"3727",x"0002",x"4784",x"4A1D",x"A003",x"FFFA",x"372A",x"0005", -- 11F0-11FF 
  x"4784",x"49FB",x"A003",x"FFFA",x"3730",x"0004",x"4784",x"4A25",x"A003",x"FFFA",x"3735",x"0001",x"4784",x"4F1F",x"A003",x"FFFA", -- 1200-120F 
  x"3737",x"0001",x"4784",x"4BE1",x"A003",x"FFFA",x"3739",x"0001",x"4784",x"4BE9",x"A003",x"FFFA",x"373B",x"0001",x"4784",x"4BF0", -- 1210-121F 
  x"A003",x"FFFA",x"373D",x"0001",x"4784",x"4D0E",x"A003",x"FFFA",x"373F",x"0004",x"4784",x"4C02",x"47A4",x"47A4",x"4A25",x"4D1C", -- 1220-122F 
  x"A003",x"FFF6",x"3744",x"0003",x"4784",x"4D29",x"A003",x"FFFA",x"3748",x"0002",x"4784",x"4D3B",x"A003",x"FFFA",x"374B",x"0001", -- 1230-123F 
  x"4784",x"4DE3",x"A003",x"FFFA",x"374D",x"0001",x"4784",x"A00A",x"520D",x"A003",x"A003",x"FFFA",x"374D",x"0001",x"478C",x"A00A", -- 1240-124F 
  SHA(10*16-1 downto 9*16),
  SHA(9*16-1 downto 8*16),
  SHA(8*16-1 downto 7*16),
  SHA(7*16-1 downto 6*16),
  SHA(6*16-1 downto 5*16),
  SHA(5*16-1 downto 4*16),
  SHA(4*16-1 downto 3*16),
  SHA(3*16-1 downto 2*16),
  SHA(2*16-1 downto 1*16),
  SHA(1*16-1 downto 0*16),
  others=>x"0000");

-- Textspeicher
type ByteRAMTYPE is array(0 to 4*1024-1) of STD_LOGIC_VECTOR (7 downto 0);
signal ByteRAM: ByteRAMTYPE:=(
  x"28",x"20",x"7B",x"20",x"7D",x"20",x"43",x"4F",x"4D",x"50",x"49",x"4C",x"45",x"20",x"28",x"4C", -- 3000-300F 
  x"49",x"54",x"2C",x"29",x"20",x"4C",x"49",x"54",x"2C",x"20",x"28",x"43",x"4F",x"4E",x"53",x"54", -- 3010-301F 
  x"41",x"4E",x"54",x"3A",x"29",x"20",x"43",x"4F",x"4E",x"53",x"54",x"41",x"4E",x"54",x"20",x"4B", -- 3020-302F 
  x"45",x"59",x"41",x"44",x"52",x"20",x"53",x"50",x"20",x"52",x"50",x"20",x"50",x"43",x"20",x"58", -- 3030-303F 
  x"42",x"49",x"54",x"20",x"53",x"4D",x"55",x"44",x"47",x"45",x"42",x"49",x"54",x"20",x"52",x"50", -- 3040-304F 
  x"30",x"20",x"49",x"52",x"41",x"4D",x"41",x"44",x"52",x"20",x"4A",x"52",x"41",x"4D",x"41",x"44", -- 3050-305F 
  x"52",x"20",x"58",x"4F",x"46",x"46",x"20",x"43",x"52",x"42",x"5A",x"45",x"49",x"47",x"20",x"43", -- 3060-306F 
  x"52",x"44",x"50",x"20",x"42",x"41",x"53",x"45",x"20",x"54",x"49",x"42",x"20",x"49",x"4E",x"31", -- 3070-307F 
  x"20",x"49",x"4E",x"32",x"20",x"49",x"4E",x"33",x"20",x"49",x"4E",x"34",x"20",x"45",x"52",x"52", -- 3080-308F 
  x"4F",x"52",x"4E",x"52",x"20",x"44",x"50",x"20",x"53",x"54",x"41",x"54",x"20",x"4C",x"46",x"41", -- 3090-309F 
  x"20",x"42",x"41",x"4E",x"46",x"20",x"42",x"5A",x"45",x"49",x"47",x"20",x"44",x"50",x"4D",x"45", -- 30A0-30AF 
  x"52",x"4B",x"20",x"43",x"53",x"50",x"20",x"44",x"55",x"42",x"49",x"54",x"20",x"4C",x"4F",x"43", -- 30B0-30BF 
  x"41",x"4C",x"41",x"44",x"52",x"45",x"53",x"53",x"45",x"20",x"56",x"45",x"52",x"53",x"49",x"4F", -- 30C0-30CF 
  x"4E",x"20",x"52",x"45",x"54",x"55",x"52",x"4E",x"20",x"28",x"4D",x"43",x"4F",x"44",x"45",x"3A", -- 30D0-30DF 
  x"29",x"20",x"4D",x"43",x"4F",x"44",x"45",x"20",x"4D",x"49",x"4E",x"55",x"53",x"20",x"55",x"2B", -- 30E0-30EF 
  x"20",x"55",x"2A",x"20",x"30",x"3D",x"20",x"30",x"4C",x"54",x"20",x"45",x"4D",x"49",x"54",x"43", -- 30F0-30FF 
  x"4F",x"44",x"45",x"20",x"4E",x"4F",x"54",x"20",x"41",x"4E",x"44",x"20",x"4F",x"52",x"20",x"2B", -- 3100-310F 
  x"20",x"21",x"20",x"40",x"20",x"53",x"57",x"41",x"50",x"20",x"4F",x"56",x"45",x"52",x"20",x"44", -- 3110-311F 
  x"55",x"50",x"20",x"52",x"4F",x"54",x"20",x"44",x"52",x"4F",x"50",x"20",x"32",x"53",x"57",x"41", -- 3120-312F 
  x"50",x"20",x"32",x"4F",x"56",x"45",x"52",x"20",x"32",x"44",x"55",x"50",x"20",x"32",x"44",x"52", -- 3130-313F 
  x"4F",x"50",x"20",x"4E",x"4F",x"4F",x"50",x"20",x"42",x"2C",x"20",x"5A",x"2C",x"20",x"28",x"57", -- 3140-314F 
  x"4F",x"52",x"44",x"3A",x"29",x"20",x"57",x"4F",x"52",x"44",x"3A",x"20",x"22",x"20",x"2E",x"22", -- 3150-315F 
  x"20",x"48",x"45",x"52",x"45",x"20",x"4A",x"52",x"42",x"49",x"54",x"20",x"4A",x"52",x"30",x"42", -- 3160-316F 
  x"49",x"54",x"20",x"58",x"53",x"45",x"54",x"42",x"54",x"20",x"41",x"4C",x"4C",x"4F",x"54",x"20", -- 3170-317F 
  x"42",x"52",x"41",x"4E",x"43",x"48",x"2C",x"20",x"30",x"42",x"52",x"41",x"4E",x"43",x"48",x"2C", -- 3180-318F 
  x"20",x"42",x"45",x"47",x"49",x"4E",x"20",x"41",x"47",x"41",x"49",x"4E",x"20",x"55",x"4E",x"54", -- 3190-319F 
  x"49",x"4C",x"20",x"49",x"46",x"20",x"45",x"4E",x"44",x"5F",x"49",x"46",x"20",x"45",x"4C",x"53", -- 31A0-31AF 
  x"45",x"20",x"57",x"48",x"49",x"4C",x"45",x"20",x"52",x"45",x"50",x"45",x"41",x"54",x"20",x"43", -- 31B0-31BF 
  x"40",x"20",x"43",x"21",x"20",x"31",x"2B",x"20",x"2D",x"20",x"3D",x"20",x"4C",x"54",x"20",x"3E", -- 31C0-31CF 
  x"20",x"2A",x"20",x"42",x"59",x"45",x"20",x"42",x"59",x"45",x"20",x"20",x"2B",x"21",x"20",x"52", -- 31D0-31DF 
  x"3E",x"20",x"3E",x"52",x"20",x"52",x"20",x"2C",x"20",x"45",x"58",x"45",x"43",x"55",x"54",x"45", -- 31E0-31EF 
  x"20",x"4B",x"45",x"59",x"20",x"45",x"4D",x"49",x"54",x"20",x"53",x"48",x"4C",x"31",x"36",x"20", -- 31F0-31FF 
  x"44",x"49",x"47",x"20",x"54",x"59",x"50",x"45",x"20",x"48",x"47",x"2E",x"20",x"48",x"2E",x"20", -- 3200-320F 
  x"2E",x"20",x"3F",x"20",x"43",x"52",x"20",x"66",x"6C",x"3E",x"20",x"2F",x"66",x"6C",x"3E",x"20", -- 3210-321F 
  x"66",x"72",x"3E",x"20",x"2F",x"66",x"72",x"3E",x"20",x"46",x"45",x"48",x"4C",x"45",x"52",x"54", -- 3220-322F 
  x"45",x"58",x"54",x"20",x"44",x"49",x"53",x"41",x"42",x"4C",x"45",x"20",x"77",x"65",x"69",x"74", -- 3230-323F 
  x"65",x"72",x"20",x"6E",x"61",x"63",x"68",x"20",x"54",x"61",x"73",x"74",x"65",x"20",x"45",x"53", -- 3240-324F 
  x"43",x"41",x"50",x"45",x"20",x"20",x"45",x"52",x"52",x"4F",x"52",x"20",x"3F",x"3F",x"3F",x"20", -- 3250-325F 
  x"46",x"45",x"48",x"4C",x"45",x"52",x"54",x"45",x"58",x"54",x"20",x"45",x"52",x"52",x"4F",x"52", -- 3260-326F 
  x"20",x"2D",x"20",x"46",x"65",x"68",x"6C",x"65",x"72",x"20",x"4E",x"75",x"6D",x"6D",x"65",x"72", -- 3270-327F 
  x"20",x"20",x"43",x"53",x"50",x"21",x"20",x"43",x"53",x"50",x"3F",x"20",x"4C",x"4F",x"43",x"41", -- 3280-328F 
  x"4C",x"20",x"45",x"4E",x"44",x"5F",x"4C",x"4F",x"43",x"41",x"4C",x"20",x"4C",x"30",x"20",x"4C", -- 3290-329F 
  x"31",x"20",x"4C",x"32",x"20",x"4C",x"33",x"20",x"4C",x"34",x"20",x"4C",x"35",x"20",x"4C",x"36", -- 32A0-32AF 
  x"20",x"4C",x"37",x"20",x"27",x"20",x"49",x"4E",x"43",x"52",x"34",x"20",x"4B",x"45",x"59",x"5F", -- 32B0-32BF 
  x"49",x"4E",x"54",x"20",x"4B",x"45",x"59",x"43",x"4F",x"44",x"45",x"32",x"20",x"45",x"58",x"50", -- 32C0-32CF 
  x"45",x"43",x"54",x"20",x"44",x"49",x"47",x"49",x"54",x"20",x"4E",x"55",x"4D",x"42",x"45",x"52", -- 32D0-32DF 
  x"20",x"57",x"4F",x"52",x"44",x"20",x"5A",x"3D",x"20",x"46",x"49",x"4E",x"44",x"20",x"4C",x"43", -- 32E0-32EF 
  x"46",x"41",x"20",x"43",x"4F",x"4D",x"50",x"49",x"4C",x"45",x"2C",x"20",x"43",x"52",x"45",x"41", -- 32F0-32FF 
  x"54",x"45",x"20",x"49",x"4E",x"54",x"45",x"52",x"50",x"52",x"45",x"54",x"20",x"51",x"55",x"49", -- 3300-330F 
  x"54",x"20",x"2F",x"6F",x"6B",x"3E",x"20",x"6F",x"6B",x"20",x"6F",x"6B",x"3E",x"20",x"2F",x"6F", -- 3310-331F 
  x"6B",x"3E",x"20",x"6F",x"6B",x"20",x"53",x"54",x"41",x"52",x"54",x"20",x"46",x"4F",x"52",x"54", -- 3320-332F 
  x"59",x"2D",x"46",x"4F",x"52",x"54",x"48",x"20",x"53",x"4D",x"55",x"44",x"47",x"45",x"20",x"28", -- 3330-333F 
  x"49",x"4D",x"4D",x"45",x"44",x"49",x"41",x"54",x"45",x"3A",x"29",x"20",x"28",x"43",x"4F",x"4D", -- 3340-334F 
  x"50",x"49",x"4C",x"45",x"3A",x"29",x"20",x"28",x"3A",x"29",x"20",x"49",x"4D",x"4D",x"45",x"44", -- 3350-335F 
  x"49",x"41",x"54",x"45",x"3A",x"20",x"43",x"4F",x"4D",x"50",x"49",x"4C",x"45",x"3A",x"20",x"3A", -- 3360-336F 
  x"20",x"3B",x"20",x"4C",x"47",x"2E",x"20",x"4E",x"47",x"2E",x"20",x"78",x"20",x"2C",x"20",x"44", -- 3370-337F 
  x"55",x"4D",x"50",x"5A",x"20",x"27",x"20",x"53",x"54",x"41",x"52",x"54",x"20",x"20",x"44",x"55", -- 3380-338F 
  x"4D",x"50",x"5A",x"3E",x"20",x"20",x"20",x"20",x"20",x"2D",x"2D",x"20",x"20",x"2D",x"20",x"2F", -- 3390-339F 
  x"44",x"55",x"4D",x"50",x"5A",x"3E",x"20",x"52",x"41",x"4D",x"50",x"31",x"20",x"56",x"41",x"52", -- 33A0-33AF 
  x"49",x"41",x"42",x"4C",x"45",x"20",x"4D",x"4F",x"56",x"45",x"20",x"46",x"49",x"4C",x"4C",x"20", -- 33B0-33BF 
  x"44",x"55",x"4D",x"50",x"20",x"4D",x"41",x"58",x"20",x"4D",x"49",x"4E",x"20",x"41",x"42",x"53", -- 33C0-33CF 
  x"20",x"4D",x"55",x"4C",x"54",x"5F",x"49",x"20",x"4D",x"55",x"4C",x"54",x"5F",x"49",x"49",x"20", -- 33D0-33DF 
  x"53",x"55",x"50",x"45",x"52",x"4D",x"55",x"4C",x"54",x"20",x"41",x"20",x"42",x"20",x"43",x"20", -- 33E0-33EF 
  x"53",x"4D",x"55",x"4C",x"20",x"41",x"44",x"44",x"49",x"45",x"52",x"20",x"44",x"49",x"33",x"32", -- 33F0-33FF 
  x"20",x"44",x"49",x"56",x"33",x"32",x"20",x"2F",x"4D",x"4F",x"44",x"20",x"2F",x"4D",x"4F",x"44", -- 3400-340F 
  x"20",x"2F",x"20",x"4D",x"4F",x"44",x"20",x"53",x"44",x"49",x"56",x"20",x"4F",x"50",x"45",x"52", -- 3410-341F 
  x"41",x"4E",x"44",x"31",x"20",x"4F",x"50",x"45",x"52",x"41",x"4E",x"44",x"32",x"20",x"45",x"52", -- 3420-342F 
  x"47",x"45",x"42",x"4E",x"49",x"53",x"20",x"5A",x"41",x"48",x"4C",x"45",x"4E",x"53",x"50",x"45", -- 3430-343F 
  x"49",x"43",x"48",x"45",x"52",x"20",x"53",x"50",x"45",x"49",x"43",x"48",x"45",x"52",x"45",x"4E", -- 3440-344F 
  x"44",x"45",x"20",x"53",x"43",x"48",x"49",x"45",x"42",x"20",x"53",x"4C",x"58",x"2D",x"3E",x"45", -- 3450-345F 
  x"52",x"47",x"45",x"42",x"4E",x"49",x"53",x"20",x"4F",x"50",x"45",x"52",x"41",x"4E",x"44",x"2D", -- 3460-346F 
  x"3E",x"53",x"4C",x"58",x"20",x"53",x"50",x"45",x"49",x"43",x"48",x"45",x"52",x"48",x"4F",x"4C", -- 3470-347F 
  x"20",x"32",x"4F",x"50",x"45",x"52",x"41",x"4E",x"44",x"45",x"4E",x"2D",x"3E",x"32",x"53",x"4C", -- 3480-348F 
  x"58",x"20",x"4E",x"2B",x"20",x"4E",x"2D",x"20",x"4E",x"2A",x"20",x"52",x"45",x"43",x"55",x"52", -- 3490-349F 
  x"53",x"45",x"20",x"4E",x"2F",x"4D",x"4F",x"44",x"20",x"48",x"47",x"30",x"2E",x"20",x"4E",x"2E", -- 34A0-34AF 
  x"20",x"2D",x"20",x"4E",x"42",x"2E",x"20",x"42",x"4C",x"4F",x"43",x"4B",x"41",x"4E",x"46",x"41", -- 34B0-34BF 
  x"4E",x"47",x"20",x"42",x"4C",x"4F",x"43",x"4B",x"45",x"4E",x"44",x"45",x"20",x"4E",x"45",x"42", -- 34C0-34CF 
  x"45",x"4E",x"52",x"45",x"43",x"48",x"4E",x"55",x"4E",x"47",x"20",x"48",x"41",x"55",x"50",x"54", -- 34D0-34DF 
  x"52",x"45",x"43",x"48",x"4E",x"55",x"4E",x"47",x"20",x"52",x"45",x"43",x"48",x"45",x"4E",x"42", -- 34E0-34EF 
  x"4C",x"4F",x"43",x"4B",x"20",x"49",x"4E",x"49",x"54",x"20",x"41",x"2B",x"30",x"20",x"42",x"2B", -- 34F0-34FF 
  x"30",x"20",x"4E",x"2F",x"20",x"4E",x"4D",x"4F",x"44",x"20",x"4E",x"47",x"47",x"54",x"20",x"4E", -- 3500-350F 
  x"42",x"4B",x"20",x"4E",x"4E",x"55",x"4D",x"42",x"45",x"52",x"20",x"4E",x"22",x"20",x"4E",x"5E", -- 3510-351F 
  x"20",x"4E",x"2E",x"20",x"2D",x"20",x"30",x"20",x"20",x"4E",x"42",x"2E",x"20",x"5A",x"45",x"52", -- 3520-352F 
  x"4C",x"45",x"47",x"20",x"4F",x"42",x"4A",x"3F",x"20",x"4C",x"20",x"47",x"20",x"48",x"20",x"4F", -- 3530-353F 
  x"2E",x"20",x"5B",x"20",x"20",x"5D",x"20",x"20",x"53",x"50",x"4D",x"45",x"52",x"4B",x"20",x"5B", -- 3540-354F 
  x"20",x"5D",x"20",x"4F",x"42",x"4A",x"2B",x"30",x"20",x"4F",x"42",x"4A",x"44",x"55",x"4D",x"50", -- 3550-355F 
  x"20",x"49",x"4E",x"56",x"45",x"52",x"54",x"49",x"45",x"52",x"45",x"4E",x"20",x"56",x"41",x"4E", -- 3560-356F 
  x"44",x"45",x"52",x"4D",x"4F",x"4E",x"44",x"45",x"4D",x"41",x"54",x"52",x"49",x"58",x"20",x"56", -- 3570-357F 
  x"4C",x"49",x"53",x"54",x"20",x"57",x"4C",x"49",x"53",x"54",x"20",x"52",x"45",x"54",x"55",x"52", -- 3580-358F 
  x"4E",x"20",x"52",x"45",x"50",x"4C",x"41",x"43",x"45",x"3A",x"20",x"46",x"4F",x"52",x"47",x"45", -- 3590-359F 
  x"54",x"20",x"6E",x"69",x"63",x"68",x"74",x"20",x"67",x"65",x"66",x"75",x"6E",x"64",x"65",x"6E", -- 35A0-35AF 
  x"20",x"20",x"46",x"45",x"48",x"4C",x"45",x"52",x"54",x"45",x"58",x"54",x"20",x"44",x"69",x"76", -- 35B0-35BF 
  x"69",x"73",x"69",x"6F",x"6E",x"20",x"64",x"75",x"72",x"63",x"68",x"20",x"4E",x"75",x"6C",x"6C", -- 35C0-35CF 
  x"20",x"57",x"6F",x"72",x"74",x"20",x"6E",x"69",x"63",x"68",x"74",x"20",x"64",x"65",x"66",x"69", -- 35D0-35DF 
  x"6E",x"69",x"65",x"72",x"74",x"20",x"45",x"69",x"6E",x"67",x"61",x"62",x"65",x"7A",x"65",x"69", -- 35E0-35EF 
  x"6C",x"65",x"20",x"7A",x"75",x"20",x"6C",x"61",x"6E",x"67",x"20",x"53",x"74",x"72",x"75",x"6B", -- 35F0-35FF 
  x"74",x"75",x"72",x"66",x"65",x"68",x"6C",x"65",x"72",x"20",x"69",x"6E",x"20",x"49",x"46",x"20", -- 3600-360F 
  x"45",x"4E",x"44",x"5F",x"49",x"46",x"20",x"42",x"45",x"47",x"49",x"4E",x"20",x"55",x"4E",x"54", -- 3610-361F 
  x"49",x"4C",x"20",x"44",x"4F",x"20",x"4C",x"4F",x"4F",x"50",x"20",x"20",x"6E",x"65",x"67",x"61", -- 3620-362F 
  x"74",x"69",x"76",x"65",x"72",x"20",x"45",x"78",x"70",x"6F",x"6E",x"65",x"6E",x"74",x"20",x"5A", -- 3630-363F 
  x"61",x"68",x"6C",x"65",x"6E",x"73",x"70",x"65",x"69",x"63",x"68",x"65",x"72",x"20",x"76",x"6F", -- 3640-364F 
  x"6C",x"6C",x"20",x"67",x"72",x"6F",x"C3",x"9F",x"65",x"20",x"67",x"61",x"6E",x"7A",x"65",x"20", -- 3650-365F 
  x"5A",x"61",x"68",x"6C",x"65",x"6E",x"20",x"6B",x"6F",x"6D",x"70",x"69",x"6C",x"69",x"65",x"72", -- 3660-366F 
  x"65",x"6E",x"20",x"67",x"65",x"68",x"74",x"20",x"6D",x"6F",x"6D",x"65",x"6E",x"74",x"61",x"6E", -- 3670-367F 
  x"20",x"6E",x"69",x"63",x"68",x"74",x"2C",x"20",x"73",x"69",x"65",x"68",x"65",x"20",x"54",x"45", -- 3680-368F 
  x"53",x"54",x"46",x"55",x"45",x"52",x"4E",x"45",x"55",x"45",x"53",x"2E",x"54",x"58",x"54",x"20", -- 3690-369F 
  x"53",x"54",x"52",x"47",x"3A",x"20",x"5E",x"47",x"20",x"2F",x"31",x"78",x"50",x"49",x"45",x"50", -- 36A0-36AF 
  x"2F",x"20",x"5E",x"46",x"20",x"51",x"55",x"49",x"54",x"20",x"5E",x"41",x"20",x"41",x"6E",x"67", -- 36B0-36BF 
  x"65",x"68",x"61",x"6C",x"74",x"65",x"6E",x"20",x"66",x"C3",x"BC",x"72",x"20",x"67",x"65",x"6E", -- 36C0-36CF 
  x"61",x"75",x"20",x"65",x"69",x"6E",x"65",x"20",x"45",x"69",x"6E",x"67",x"61",x"62",x"65",x"7A", -- 36D0-36DF 
  x"65",x"69",x"6C",x"65",x"3A",x"20",x"20",x"6F",x"6B",x"20",x"51",x"55",x"45",x"52",x"59",x"20", -- 36E0-36EF 
  x"28",x"2A",x"52",x"45",x"4D",x"2A",x"29",x"20",x"2F",x"6F",x"6B",x"3E",x"20",x"28",x"2A",x"45", -- 36F0-36FF 
  x"4E",x"44",x"2A",x"29",x"20",x"6F",x"6B",x"3E",x"20",x"48",x"45",x"58",x"20",x"44",x"45",x"43", -- 3700-370F 
  x"49",x"4D",x"41",x"4C",x"20",x"4E",x"4C",x"49",x"54",x"2C",x"20",x"4D",x"2E",x"20",x"4D",x"2B", -- 3710-371F 
  x"20",x"4D",x"2D",x"20",x"4D",x"2A",x"20",x"4D",x"2F",x"20",x"4D",x"2F",x"4D",x"4F",x"44",x"20", -- 3720-372F 
  x"4D",x"4D",x"4F",x"44",x"20",x"2E",x"20",x"2B",x"20",x"2D",x"20",x"2A",x"20",x"2F",x"20",x"2F", -- 3730-373F 
  x"4D",x"4F",x"44",x"20",x"47",x"47",x"54",x"20",x"42",x"4B",x"20",x"5E",x"20",x"3F",x"20",x"4D", -- 3740-374F 
  others=>x"00");

-- Rückkehrstapel
type stapRAMTYPE is array(0 to 1024-1) of STD_LOGIC_VECTOR (15 downto 0);
shared variable stapR: stapRAMTYPE:=(
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C00-2C0F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C10-2C1F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C20-2C2F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C30-2C3F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C40-2C4F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C50-2C5F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C60-2C6F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C70-2C7F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C80-2C8F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C90-2C9F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2CA0-2CAF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2CB0-2CBF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2CC0-2CCF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2CD0-2CDF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2CE0-2CEF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2CF0-2CFF 
  x"0000",x"0000",x"0000",x"0000",x"0055",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D00-2D0F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D10-2D1F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D20-2D2F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D30-2D3F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D40-2D4F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D50-2D5F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D60-2D6F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D70-2D7F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D80-2D8F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D90-2D9F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2DA0-2DAF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2DB0-2DBF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2DC0-2DCF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2DD0-2DDF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2DE0-2DEF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2DF0-2DFF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E00-2E0F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E10-2E1F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E20-2E2F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E30-2E3F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E40-2E4F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E50-2E5F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E60-2E6F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E70-2E7F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E80-2E8F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E90-2E9F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2EA0-2EAF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2EB0-2EBF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2EC0-2ECF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2ED0-2EDF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0008", -- 2EE0-2EEF 
  x"0008",x"0000",x"0001",x"2F22",x"0000",x"0001",x"2F23",x"1410",x"0008",x"3B0A",x"0001",x"0001",x"3B45",x"00BB",x"0001",x"FFFF", -- 2EF0-2EFF 
  x"0000",x"0000",x"3000",x"3D49",x"3D49",x"FFFF",x"374F",x"124A",x"0010",x"3B00",x"3B00",x"3B0C",x"3B12",x"3B45",x"0000",x"124A", -- 2F00-2F0F 
  x"0000",x"1243",x"3000",x"374F",x"0020",x"0065",x"0000",x"2F00",x"0000",x"1190",x"0000",x"0000",x"0000",x"0000",x"1185",x"117B", -- 2F10-2F1F 
  x"2F2A",x"0000",x"0000",x"140C",x"1400",x"2000",x"0001",x"1400",x"1400",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F20-2F2F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F30-2F3F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F40-2F4F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F50-2F5F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F60-2F6F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F70-2F7F 
  x"2F00",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F80-2F8F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F90-2F9F 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2FA0-2FAF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2FB0-2FBF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2FC0-2FCF 
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0301",x"0301",x"0301",x"0301",x"0301",x"0301",x"0301",x"0301", -- 2FD0-2FDF 
  x"0301",x"0301",x"0301",x"0301",x"0446",x"02D5",x"02CD",x"004B",x"02CD",x"02CD",x"02CD",x"02CD",x"02CD",x"0655",x"02CD",x"004B", -- 2FE0-2FEF 
  x"02CD",x"02CD",x"02CD",x"004B",x"0318",x"033F",x"01EC",x"0288",x"080C",x"FFFF",x"06F1",x"3B05",x"3B06",x"3B00",x"3B00",x"073B", -- 2FF0-2FFF 
  others=>x"0000");

--diese Funktion übernimmt von SP nur die beiden niedrigsten Bits
  function P(SP : integer) return integer is begin
--    return CONV_INTEGER(CONV_UNSIGNED(SP,2));
    return SP mod 4;
    end;

-- alles Signale um die Stapel-RAM's zu machen.
signal HOLE_VOM_STAPEL,STORE_ZUM_STAPEL,ADRESSE_ZUM_STAPEL: REG;
signal WE_ZUM_STAPEL: STD_LOGIC_VECTOR (3 downto 0);
type STAPELTYPE is array(0 to 31) of STD_LOGIC_VECTOR (15 downto 0);
signal stap1,stap2,stap3,stap0: STAPELTYPE:=(others=>x"0000");
-- Rueckkehrstapel
signal RPC,RPCC: STD_LOGIC_VECTOR (15 downto 0);
signal RP: STD_LOGIC_VECTOR (15 downto 0):=x"3000";
signal RW: STD_LOGIC;
-- kompletten Speicher anschliessen
signal PC_ZUM_ProgRAM,PD_VOM_ProgRAM: STD_LOGIC_VECTOR (15 downto 0);
signal STORE_ZUM_RAM,EXFET,ADRESSE_ZUM_RAM: STD_LOGIC_VECTOR (15 downto 0);
signal FETCH_VOM_ProgRAM,FETCH_VOM_ByteRAM,FETCH_VOM_stapR: STD_LOGIC_VECTOR (15 downto 0);
signal WE_ZUM_RAM,WE_ZUM_ProgRAM,WE_ZUM_ByteRAM,WE_ZUM_stapR: STD_LOGIC;
-- fuer EMIT-Ausgabe
signal EMIT_ABGESCHICKT_LOCAL,EMIT_ANGEKOMMEN_RUHEND,XOFF_INPUT_L: STD_LOGIC:='0';
signal KEY_ANGEKOMMEN_LOCAL,KEY_ABGESCHICKT_RUHEND,KEY_ABGESCHICKT_MERK: STD_LOGIC:='0';
signal KEY_BYTE_RUHEND: STD_LOGIC_VECTOR (7 downto 0);


begin

process begin wait until (CLK_I'event and CLK_I='1'); --ruhende Eingangsdaten für FortyForthprocessor
  EMIT_ANGEKOMMEN_RUHEND<=EMIT_ANGEKOMMEN;
  KEY_BYTE_RUHEND<=KEY_BYTE;
  KEY_ABGESCHICKT_RUHEND<=KEY_ABGESCHICKT;
  end process;
  

process -- FortyForthProcessor
variable PC,PD,ADR,DAT,DIST: STD_LOGIC_VECTOR (15 downto 0):=x"0000";
variable WE: STD_LOGIC;
variable SP: integer:=0;
variable R: REG:=(others=>x"0000");
-- Stapeleintraege benennen
variable A,B,C,D: STD_LOGIC_VECTOR (15 downto 0):=x"0000";
variable T: integer range 0 to 4;
variable W: STD_LOGIC_VECTOR (3 downto 0);
-- fuer Umstapeln 
variable STAK: STD_LOGIC_VECTOR (7 downto 0);
-- fuer Rechenoperationen mit Uebertrag
variable U: STD_LOGIC_VECTOR (31 downto 0);
-- fuer Division
variable UBIT: STD_LOGIC;
-- fuer Supermult
variable SUMME: STD_LOGIC_VECTOR (31 downto 0);

begin wait until (CLK_I'event and CLK_I='0'); PC_SIM<=PC;--Simulation
  -- ob ein KEY aingetroffen ist --
  if KEY_ABGESCHICKT_MERK/=KEY_ABGESCHICKT_RUHEND then 
    KEY_ABGESCHICKT_MERK<=KEY_ABGESCHICKT_RUHEND;
    PD:=x"4012";
    PC:=PC;
    else
      PD:=PD_VOM_ProgRAM;
      PC:=PC+1;
      end if;                                           -- Simulation --
  WE:='0';                                              PD_SIM<=PD;
  DIST:=PD(11)&PD(11)&PD(11)&PD(11)&PD(11 downto 0);    SP_SIM<=SP;
  -- oberste 4 Stapeleintraege entnehmen
  R:=HOLE_VOM_STAPEL;                                   -- Simulation --
  A:=R(P(SP-1));                                        A_SIM<=A;
  B:=R(P(SP-2));                                        B_SIM<=B;
  C:=R(P(SP-3));                                        C_SIM<=C;
  D:=R(P(SP-4));                                        D_SIM<=D;
  T:=0;
  -- Rueckkehrstapel
  RW<='0';
 
  if PD(15 downto 13)="010" then                 -- 4000-5FFF Unterprogrammaufruf
    RPC<=PC;PC:=PD and x"3FFF";RP<=RP-1;RW<='1';
    elsif PD(15 downto 12)=x"8" then PC:=PC+DIST;-- 8000-8FFF relativer Sprung
    elsif PD(15 downto 12)=x"9" then             -- 9000-9FFF bedingter relativer Sprung
      if A=x"0000" then PC:=PC+DIST; end if; SP:=SP-1;
    elsif PD=x"A003" then PC:=RPCC;RP<=RP+1;     -- ; Rückkehr aus Unterprogramm
    elsif PD=x"A00D" then -- 0= Vergleich ob gleich Null
      if A=x"0000" then A:=x"FFFF"; 
        else A:=x"0000"; end if;
      T:=1;
    elsif PD=x"A00F" then -- 0< Vergleich ob kleiner Null
      if A>=x"8000" then A:=x"FFFF";
        else A:=x"0000"; end if;
      T:=1;
    elsif PD=x"A000" then -- MINUS Vorzeichen wechseln
      A:=(not A)+1;
      T:=1;
    elsif PD=x"A00B" then -- NOT Bitweises Komplement
      A:=not A;
      T:=1;
    elsif PD=x"A008" then -- AND Bitweises Und
      A:=B and A; 
      T:=1;
      SP:=SP-1;
    elsif PD=x"A00E" then -- OR Bitweises Oder
      A:=B or A; 
      T:=1;
      SP:=SP-1;
    elsif PD=x"A007" then -- + Addition
      A:=B+A; 
      T:=1;
      SP:=SP-1;
    elsif PD=x"A001" then -- U+ Addition mit Übertrag
      U:=(x"0000"&C)+(x"0000"&B)+(x"0000"&A);
      B:=U(31 downto 16);
      A:=U(15 downto 0);
      T:=2;
      SP:=SP-1;
    elsif PD=x"A002" then -- U* Multiplikation mit Übertrag
      U:=(x"0000"&C)+B*A;
      B:=U(31 downto 16);
      A:=U(15 downto 0);
      T:=2;
      SP:=SP-1;
    elsif PD=x"A005" then -- EMIT Zeichen ausgeben
      if (EMIT_ABGESCHICKT_LOCAL=EMIT_ANGEKOMMEN_RUHEND) and XOFF_INPUT_L='0' then
        EMIT_BYTE<=A(7 downto 0);
        EMIT_ABGESCHICKT_LOCAL<=not EMIT_ANGEKOMMEN_RUHEND;
        T:=0;
        SP:=SP-1;
        else PC:=PC-1; end if; -- warten
    elsif PD=x"A009" then -- STORE Speicheradresse beschreiben
      case A is
        when x"2800" => KEY_ANGEKOMMEN_LOCAL<=not KEY_ANGEKOMMEN_LOCAL;
        when x"2801" => SP:=CONV_INTEGER(B);
        when x"2802" => RP<=B;
        when x"2803" => PC:=B;
        when others => ADR:=A;DAT:=B;WE:='1' ;
        end case;
      T:=0;
      SP:=SP-2;
    elsif PD=x"A00A" then -- FETCH Speicheradresse lesen
      case A is
        when x"2800" => A:=x"00"&KEY_BYTE_RUHEND;
        when x"2801" => A:=CONV_STD_LOGIC_VECTOR(SP-1,16);
        when x"2802" => A:=RP;
        when x"2803" => A:=PC;
        when others => A:=EXFET;
        end case;
      T:=1;
    elsif PD=x"A014" then -- DI32 DIVISION_MIT_REST 32B/16B=16R/16Q
      UBIT:=C(15);
      C:=C(14 downto 0)&B(15);
      B:=B(14 downto 0)&'0';
      if (UBIT&C)>=('0'&A) then
        C:=C-A;
        B(0):='1';
        end if;
      T:=3;
    elsif PD=x"A017" then -- MULT_I
      --     D    C    B    A        stapR
      --     c    ü   adr1 adr2      i
      -- c   ü   erg1 adr2 adr1      i-1
      SUMME:=(D*EXFET)+(x"0000"&C);
      C:=A;A:=B;B:=C;
      D:=SUMME(31 downto 16); 
      C:=SUMME(15 downto 0);
      RPC<=RPCC-1; RW<='1';
      T:=4; SP:=SP+1;
    elsif PD=x"A018" then -- MULT_II
      --     D    C     B      A         stapR
      -- c   ü1  erg1   adr2   adr1      i-1
      -- c   ü2  adr1+1 adr2+1 i-1       i-1
      SUMME:=(D&C)+(x"0000"&EXFET);
      D:=SUMME(31 downto 16); 
      DAT:=SUMME(15 downto 0);
      ADR:=A;
      WE:='1';
      C:=A+1;
      B:=B+1;
      if RPCC=x"0000" then A:=x"FFFF"; else A:=x"0000"; end if;
      T:=4;
    elsif PD(15 downto 12)=x"B" then           -- B000-BFFF Umstapeln
      STAK:="00000000";
      if PD(7)='1' then STAK:=STAK(5 downto 0)&"11"; T:=T+1; end if;
      if PD(6)='1' then STAK:=STAK(5 downto 0)&"10"; T:=T+1; end if;
      if PD(5)='1' then STAK:=STAK(5 downto 0)&"01"; T:=T+1; end if;
      if PD(4)='1' then STAK:=STAK(5 downto 0)&"00"; T:=T+1; end if;
      if PD(3)='1' then STAK:=STAK(5 downto 0)&"11"; T:=T+1; end if;
      if PD(2)='1' then STAK:=STAK(5 downto 0)&"10"; T:=T+1; end if;
      if PD(1)='1' then STAK:=STAK(5 downto 0)&"01"; T:=T+1; end if;
      if PD(0)='1' then STAK:=STAK(5 downto 0)&"00"; T:=T+1; end if;
      A:=R(P(SP-1-CONV_INTEGER(STAK(1 downto 0))));
      B:=R(P(SP-1-CONV_INTEGER(STAK(3 downto 2))));
      C:=R(P(SP-1-CONV_INTEGER(STAK(5 downto 4))));
      D:=R(P(SP-1-CONV_INTEGER(STAK(7 downto 6))));
      SP:=SP+CONV_INTEGER(PD(11 downto 8))-4;
    else A:=PD; SP:=SP+1; T:=1; end if;                    -- LIT
    
  -- oberste T Stapeleintraege zurückspeichern
  W:="0000";
  if T/=0 then R(P(SP-1)):=A; W(P(SP-1)):='1';
    if T/=1 then R(P(SP-2)):=B; W(P(SP-2)):='1';
      if T/=2 then R(P(SP-3)):=C; W(P(SP-3)):='1';
        if T/=3 then R(P(SP-4)):=D; W(P(SP-4)):='1';
          end if; end if; end if; end if;
  -- Ausgabeadresse zum StapRAM zusammenbasteln
  ADRESSE_ZUM_STAPEL(0)<=CONV_STD_LOGIC_VECTOR(SP-1,16);
  ADRESSE_ZUM_STAPEL(1)<=CONV_STD_LOGIC_VECTOR(SP-2,16);
  ADRESSE_ZUM_STAPEL(2)<=CONV_STD_LOGIC_VECTOR(SP-3,16);
  ADRESSE_ZUM_STAPEL(3)<=CONV_STD_LOGIC_VECTOR(SP-4,16);
  STORE_ZUM_STAPEL<=R;
  WE_ZUM_STAPEL<=W;
  -- ADR, DAT, WE, PC
  if WE='1' then ADRESSE_ZUM_RAM<=ADR; else ADRESSE_ZUM_RAM<=R(P(SP-1)); end if;
  STORE_ZUM_RAM<=DAT;
  WE_ZUM_RAM<=WE;
  PC_ZUM_ProgRAM<=PC;
  end process;

ADR_O<=ADRESSE_ZUM_RAM;
DAT_O<=STORE_ZUM_RAM;
WE_O<=WE_ZUM_RAM;
EMIT_ABGESCHICKT<=EMIT_ABGESCHICKT_LOCAL;
KEY_ANGEKOMMEN<=KEY_ANGEKOMMEN_LOCAL;

-- hier werden die Lesedaten der unterschiedlichen Speicher zusammengefuehrt
EXFET<=FETCH_VOM_ProgRAM when ADRESSE_ZUM_RAM(15 downto 13)="000" else
       FETCH_VOM_stapR when ADRESSE_ZUM_RAM(15 downto 10)="001011" else
       x"00"&FETCH_VOM_ByteRAM(7 downto 0) when ADRESSE_ZUM_RAM(15 downto 12)="0011" else
       DAT_I;

-- hier wird WE auf die unterschiedlichen Speicher aufgeteilt
WE_ZUM_ProgRAM<=WE_ZUM_RAM when ADRESSE_ZUM_RAM(15 downto 13)="000" else '0';
WE_ZUM_stapR  <=WE_ZUM_RAM when ADRESSE_ZUM_RAM(15 downto 10)="001011" else '0';
WE_ZUM_ByteRAM<=WE_ZUM_RAM when ADRESSE_ZUM_RAM(15 downto 12)="0011" else '0';


process -- Programmspeicher 0000H-1FFFH,
begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_ProgRAM='1' then 
    ProgRAM(CONV_INTEGER(ADRESSE_ZUM_RAM(12 downto 0)))<=STORE_ZUM_RAM; 
    FETCH_VOM_ProgRAM<=STORE_ZUM_RAM; 
	  else
      FETCH_VOM_ProgRAM<=ProgRAM(CONV_INTEGER(ADRESSE_ZUM_RAM(12 downto 0)));
      end if;
  PD_VOM_ProgRAM<=ProgRAM(CONV_INTEGER(PC_ZUM_ProgRAM(12 downto 0)));
  end process;

process -- Textspeicher 3000H-3FFFH
begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_ByteRAM='1' then 
    ByteRAM(CONV_INTEGER(ADRESSE_ZUM_RAM(11 downto 0)))<=STORE_ZUM_RAM(7 downto 0); 
    FETCH_VOM_ByteRAM<=STORE_ZUM_RAM; 
	 else
      FETCH_VOM_ByteRAM<=x"00"&ByteRAM(CONV_INTEGER(ADRESSE_ZUM_RAM(11 downto 0)));
      end if;
  end process;

process --Rueckkehrstapel, TRUE_DUAL_PORT
begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_StapR='1' then 
    stapR(CONV_INTEGER(ADRESSE_ZUM_RAM(9 downto 0))):=STORE_ZUM_RAM; 
    end if;
  FETCH_VOM_stapR<=stapR(CONV_INTEGER(ADRESSE_ZUM_RAM(9 downto 0)));
  end process;
process begin wait until (CLK_I'event and CLK_I='1');
  if RW='1' then
    stapR(CONV_INTEGER(RP(9 downto 0))):=RPC;
    RPCC<=RPC;
     else
      RPCC<=stapR(CONV_INTEGER(RP(9 downto 0)));
    end if;
  end process;

--StapelRAM:
process begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_STAPEL(0)='1' then
    stap0(CONV_INTEGER(ADRESSE_ZUM_STAPEL(0)(6 downto 2)))<=STORE_ZUM_STAPEL(0);
    HOLE_VOM_STAPEL(0)<=STORE_ZUM_STAPEL(0);
     else
      HOLE_VOM_STAPEL(0)<=stap0(CONV_INTEGER(ADRESSE_ZUM_STAPEL(0)(6 downto 2)));
    end if;
  end process;
process begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_STAPEL(1)='1' then
    stap1(CONV_INTEGER(ADRESSE_ZUM_STAPEL(1)(6 downto 2)))<=STORE_ZUM_STAPEL(1);
    HOLE_VOM_STAPEL(1)<=STORE_ZUM_STAPEL(1);
     else
      HOLE_VOM_STAPEL(1)<=stap1(CONV_INTEGER(ADRESSE_ZUM_STAPEL(1)(6 downto 2)));
    end if;
  end process;
process begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_STAPEL(2)='1' then
    stap2(CONV_INTEGER(ADRESSE_ZUM_STAPEL(2)(6 downto 2)))<=STORE_ZUM_STAPEL(2);
    HOLE_VOM_STAPEL(2)<=STORE_ZUM_STAPEL(2);
     else
      HOLE_VOM_STAPEL(2)<=stap2(CONV_INTEGER(ADRESSE_ZUM_STAPEL(2)(6 downto 2)));
    end if;
  end process;
process begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_STAPEL(3)='1' then
    stap3(CONV_INTEGER(ADRESSE_ZUM_STAPEL(3)(6 downto 2)))<=STORE_ZUM_STAPEL(3);
    HOLE_VOM_STAPEL(3)<=STORE_ZUM_STAPEL(3);
     else
      HOLE_VOM_STAPEL(3)<=stap3(CONV_INTEGER(ADRESSE_ZUM_STAPEL(3)(6 downto 2)));
    end if;
  end process;

end Step_9;
