library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity top is
  Port ( 
    CLK: in STD_LOGIC;
    LEDS: out STD_LOGIC_VECTOR (7 downto 0);
            
    -- EMIT --
    EMIT_ABGESCHICKT: out STD_LOGIC;
    EMIT_BYTE: out STD_LOGIC_VECTOR (7 downto 0);
    EMIT_ANGEKOMMEN: in STD_LOGIC;

     -- KEY --
    KEY_ABGESCHICKT: in STD_LOGIC;
    KEY_BYTE: in STD_LOGIC_VECTOR (7 downto 0);
    KEY_ANGEKOMMEN: out STD_LOGIC;

    -- nur zur Simulation und Fehlersuche:
    CLK_SIM : out STD_LOGIC;
    PC_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    PD_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    SP_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    A_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    B_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    C_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    D_SIM: out STD_LOGIC_VECTOR (15 downto 0)
    );
  end top;

architecture Step_1 of top is

component FortyForthProcessor
  port (
    CLK_I: in STD_LOGIC;
    DAT_I: in STD_LOGIC_VECTOR (15 downto 0);
    ADR_O: out STD_LOGIC_VECTOR (15 downto 0);
    DAT_O: out STD_LOGIC_VECTOR (15 downto 0);
    WE_O: out STD_LOGIC;
        
    -- EMIT --
    EMIT_ABGESCHICKT: out STD_LOGIC;
    EMIT_BYTE: out STD_LOGIC_VECTOR (7 downto 0);
    EMIT_ANGEKOMMEN: in STD_LOGIC;

     -- KEY --
    KEY_ABGESCHICKT: in STD_LOGIC;
    KEY_BYTE: in STD_LOGIC_VECTOR (7 downto 0);
    KEY_ANGEKOMMEN: out STD_LOGIC;

    -- LINKS --
    LINKS_ABGESCHICKT: in STD_LOGIC;
    LINKS_DAT:  in STD_LOGIC_VECTOR (15 downto 0);
    LINKS_ADR: out STD_LOGIC_VECTOR (15 downto 0);
    LINKS_ANGEKOMMEN: out STD_LOGIC;
    
    -- RECHTS --
    RECHTS_ABGESCHICKT: out STD_LOGIC;
    RECHTS_DAT: out STD_LOGIC_VECTOR (15 downto 0);
    RECHTS_ADR:  in STD_LOGIC_VECTOR (15 downto 0);
    RECHTS_ANGEKOMMEN: in STD_LOGIC;
    
    -- OBEN --
    OBEN_ABGESCHICKT: in STD_LOGIC;
    OBEN_DAT:  in STD_LOGIC_VECTOR (15 downto 0);
    OBEN_ADR: out STD_LOGIC_VECTOR (15 downto 0);
    OBEN_ANGEKOMMEN: out STD_LOGIC;
    
    -- UNTEN --
    UNTEN_ABGESCHICKT: out STD_LOGIC;
    UNTEN_DAT: out STD_LOGIC_VECTOR (15 downto 0);
    UNTEN_ADR:  in STD_LOGIC_VECTOR (15 downto 0);
    UNTEN_ANGEKOMMEN: in STD_LOGIC;
    
    -- nur zur Simulation und Fehlersuche:
    PC_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    PD_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    SP_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    A_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    B_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    C_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    D_SIM: out STD_LOGIC_VECTOR (15 downto 0)
    );
  end component;

signal WE      : STD_LOGIC;
signal ADR,DAT : STD_LOGIC_VECTOR (15 downto 0);

signal L00_AB, L00_AN, R00_AB, R00_AN, O00_AB, O00_AN, U00_AB, U00_AN:  STD_LOGIC;
signal L00_DAT,L00_ADR,R00_DAT,R00_ADR,O00_DAT,O00_ADR,U00_DAT,U00_ADR: STD_LOGIC_VECTOR (15 downto 0);
signal L01_AB, L01_AN, R01_AB, R01_AN, O01_AB, O01_AN, U01_AB, U01_AN:  STD_LOGIC;
signal L01_DAT,L01_ADR,R01_DAT,R01_ADR,O01_DAT,O01_ADR,U01_DAT,U01_ADR: STD_LOGIC_VECTOR (15 downto 0);
signal L10_AB, L10_AN, R10_AB, R10_AN, O10_AB, O10_AN, U10_AB, U10_AN:  STD_LOGIC;
signal L10_DAT,L10_ADR,R10_DAT,R10_ADR,O10_DAT,O10_ADR,U10_DAT,U10_ADR: STD_LOGIC_VECTOR (15 downto 0);
signal L11_AB, L11_AN, R11_AB, R11_AN, O11_AB, O11_AN, U11_AB, U11_AN:  STD_LOGIC;
signal L11_DAT,L11_ADR,R11_DAT,R11_ADR,O11_DAT,O11_ADR,U11_DAT,U11_ADR: STD_LOGIC_VECTOR (15 downto 0);

signal NN01,NN10,NN11: STD_LOGIC;

begin
  -- component instantiation
DUT00: FortyForthProcessor
  port map (
    CLK_I => CLK,DAT_I => x"0000",ADR_O => ADR,DAT_O => DAT,WE_O => WE,
      EMIT_ABGESCHICKT => EMIT_ABGESCHICKT,EMIT_BYTE => EMIT_BYTE,EMIT_ANGEKOMMEN => EMIT_ANGEKOMMEN,-- EMIT --
       KEY_ABGESCHICKT => KEY_ABGESCHICKT,  KEY_BYTE => KEY_BYTE,  KEY_ANGEKOMMEN => KEY_ANGEKOMMEN, -- KEY --
     LINKS_ABGESCHICKT => L00_AB, LINKS_DAT => L00_DAT, LINKS_ADR => L00_ADR, LINKS_ANGEKOMMEN => L00_AN,-- LINKS --
    RECHTS_ABGESCHICKT => R00_AB,RECHTS_DAT => R00_DAT,RECHTS_ADR => R00_ADR,RECHTS_ANGEKOMMEN => R00_AN,-- RECHTS --
      OBEN_ABGESCHICKT => O00_AB,  OBEN_DAT => O00_DAT,  OBEN_ADR => O00_ADR,  OBEN_ANGEKOMMEN => O00_AN,-- OBEN --
     UNTEN_ABGESCHICKT => U00_AB, UNTEN_DAT => U00_DAT, UNTEN_ADR => U00_ADR, UNTEN_ANGEKOMMEN => U00_AN,-- UNTEN --
    PC_SIM => PC_SIM,PD_SIM => PD_SIM,A_SIM => A_SIM,B_SIM => B_SIM,C_SIM => C_SIM,D_SIM => D_SIM,SP_SIM => SP_SIM-- nur fuer Simulation
    );

DUT01: FortyForthProcessor
  port map (
    CLK_I => CLK,DAT_I => x"0000",ADR_O => ADR,DAT_O => DAT,WE_O => WE,
      EMIT_ABGESCHICKT => NN01,EMIT_BYTE => open, EMIT_ANGEKOMMEN => NN01, -- EMIT --
       KEY_ABGESCHICKT => '0',  KEY_BYTE => x"00", KEY_ANGEKOMMEN => open, -- KEY --
     LINKS_ABGESCHICKT => L01_AB, LINKS_DAT => L01_DAT, LINKS_ADR => L01_ADR, LINKS_ANGEKOMMEN => L01_AN,-- LINKS --
    RECHTS_ABGESCHICKT => R01_AB,RECHTS_DAT => R01_DAT,RECHTS_ADR => R01_ADR,RECHTS_ANGEKOMMEN => R01_AN,-- RECHTS --
      OBEN_ABGESCHICKT => O01_AB,  OBEN_DAT => O01_DAT,  OBEN_ADR => O01_ADR,  OBEN_ANGEKOMMEN => O01_AN,-- OBEN --
     UNTEN_ABGESCHICKT => U01_AB, UNTEN_DAT => U01_DAT, UNTEN_ADR => U01_ADR, UNTEN_ANGEKOMMEN => U01_AN,-- UNTEN --
    PC_SIM =>open,PD_SIM=>open,A_SIM=>open,B_SIM=>open,C_SIM=>open,D_SIM =>open,SP_SIM=>open-- nur fuer Simulation
    );

DUT10: FortyForthProcessor
  port map (
    CLK_I => CLK,DAT_I => x"0000",ADR_O => ADR,DAT_O => DAT,WE_O => WE,
      EMIT_ABGESCHICKT => NN10,EMIT_BYTE => open, EMIT_ANGEKOMMEN => NN10, -- EMIT --
       KEY_ABGESCHICKT => '0',  KEY_BYTE => x"00", KEY_ANGEKOMMEN => open, -- KEY --
     LINKS_ABGESCHICKT => L10_AB, LINKS_DAT => L10_DAT, LINKS_ADR => L10_ADR, LINKS_ANGEKOMMEN => L10_AN,-- LINKS --
    RECHTS_ABGESCHICKT => R10_AB,RECHTS_DAT => R10_DAT,RECHTS_ADR => R10_ADR,RECHTS_ANGEKOMMEN => R10_AN,-- RECHTS --
      OBEN_ABGESCHICKT => O10_AB,  OBEN_DAT => O10_DAT,  OBEN_ADR => O10_ADR,  OBEN_ANGEKOMMEN => O10_AN,-- OBEN --
     UNTEN_ABGESCHICKT => U10_AB, UNTEN_DAT => U10_DAT, UNTEN_ADR => U10_ADR, UNTEN_ANGEKOMMEN => U10_AN,-- UNTEN --
    PC_SIM =>open,PD_SIM=>open,A_SIM=>open,B_SIM=>open,C_SIM=>open,D_SIM =>open,SP_SIM=>open-- nur fuer Simulation
    );

DUT11: FortyForthProcessor
  port map (
    CLK_I => CLK,DAT_I => x"0000",ADR_O => ADR,DAT_O => DAT,WE_O => WE,
      EMIT_ABGESCHICKT => NN11,EMIT_BYTE => open, EMIT_ANGEKOMMEN => NN11, -- EMIT --
       KEY_ABGESCHICKT => '0',  KEY_BYTE => x"00", KEY_ANGEKOMMEN => open, -- KEY --
     LINKS_ABGESCHICKT => L11_AB, LINKS_DAT => L11_DAT, LINKS_ADR => L11_ADR, LINKS_ANGEKOMMEN => L11_AN,-- LINKS --
    RECHTS_ABGESCHICKT => R11_AB,RECHTS_DAT => R11_DAT,RECHTS_ADR => R11_ADR,RECHTS_ANGEKOMMEN => R11_AN,-- RECHTS --
      OBEN_ABGESCHICKT => O11_AB,  OBEN_DAT => O11_DAT,  OBEN_ADR => O11_ADR,  OBEN_ANGEKOMMEN => O11_AN,-- OBEN --
     UNTEN_ABGESCHICKT => U11_AB, UNTEN_DAT => U11_DAT, UNTEN_ADR => U11_ADR, UNTEN_ANGEKOMMEN => U11_AN,-- UNTEN --
    PC_SIM =>open,PD_SIM=>open,A_SIM=>open,B_SIM=>open,C_SIM=>open,D_SIM =>open,SP_SIM=>open-- nur fuer Simulation
    );


L01_AB<=R00_AB; L01_DAT<=R00_DAT; R00_ADR<=L01_ADR; R00_AN<=L01_AN;
L00_AB<=R01_AB; L00_DAT<=R01_DAT; R01_ADR<=L00_ADR; R01_AN<=L00_AN;
L11_AB<=R10_AB; L11_DAT<=R10_DAT; R10_ADR<=L11_ADR; R10_AN<=L11_AN;
L10_AB<=R11_AB; L10_DAT<=R11_DAT; R11_ADR<=L10_ADR; R11_AN<=L10_AN;

O10_AB<=U00_AB; O10_DAT<=U00_DAT; O00_ADR<=U10_ADR; U00_AN<=O10_AN;
O00_AB<=U10_AB; O00_DAT<=U10_DAT; O10_ADR<=U00_ADR; U10_AN<=O00_AN;
O11_AB<=U01_AB; O11_DAT<=U01_DAT; O01_ADR<=U11_ADR; U01_AN<=O11_AN;
O01_AB<=U11_AB; O01_DAT<=U11_DAT; O11_ADR<=U01_ADR; U11_AN<=O01_AN;


process begin wait until (CLK'event and CLK='1');
  if WE='1' then
    if ADR=x"2D04" then LEDS<=DAT(7 downto 0); 
      end if; 
    end if;
  end process;

end Step_1;

