library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity FortyForthProcessor is
  Port (
    CLK_I: in STD_LOGIC;
    DAT_I: in STD_LOGIC_VECTOR (15 downto 0);
    ADR_O: out STD_LOGIC_VECTOR (15 downto 0);
    DAT_O: out STD_LOGIC_VECTOR (15 downto 0);
    WE_O: out STD_LOGIC;
    
    -- EMIT --
    EMIT_ABGESCHICKT: out STD_LOGIC;
    EMIT_BYTE: out STD_LOGIC_VECTOR (7 downto 0);
    EMIT_ANGEKOMMEN: in STD_LOGIC;
    
    -- KEY --
    KEY_ABGESCHICKT: in STD_LOGIC;
    KEY_BYTE: in STD_LOGIC_VECTOR (7 downto 0);
    KEY_ANGEKOMMEN: out STD_LOGIC;

    -- LINKS --
    LINKS_ABGESCHICKT: in STD_LOGIC;
    LINKS_DAT:  in STD_LOGIC_VECTOR (15 downto 0);
    LINKS_ADR: out STD_LOGIC_VECTOR (15 downto 0);
    LINKS_ANGEKOMMEN: out STD_LOGIC:='0';
    
    -- RECHTS --
    RECHTS_ABGESCHICKT: out STD_LOGIC:='0';
    RECHTS_DAT: out STD_LOGIC_VECTOR (15 downto 0);
    RECHTS_ADR:  in STD_LOGIC_VECTOR (15 downto 0);
    RECHTS_ANGEKOMMEN: in STD_LOGIC;
    
    -- OBEN --
    OBEN_ABGESCHICKT: in STD_LOGIC;
    OBEN_DAT:  in STD_LOGIC_VECTOR (15 downto 0);
    OBEN_ADR: out STD_LOGIC_VECTOR (15 downto 0);
    OBEN_ANGEKOMMEN: out STD_LOGIC:='0';
    
    -- UNTEN --
    UNTEN_ABGESCHICKT: out STD_LOGIC:='0';
    UNTEN_DAT: out STD_LOGIC_VECTOR (15 downto 0);
    UNTEN_ADR:  in STD_LOGIC_VECTOR (15 downto 0);
    UNTEN_ANGEKOMMEN: in STD_LOGIC;
    
   -- nur zur Simulation und Fehlersuche:
    PC_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    PD_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    SP_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    A_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    B_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    C_SIM: out STD_LOGIC_VECTOR (15 downto 0);
    D_SIM: out STD_LOGIC_VECTOR (15 downto 0)
    );
end FortyForthProcessor;

architecture Step_12 of FortyForthProcessor is

constant SHA: STD_LOGIC_VECTOR (10*16-1 downto 0):=
  x"88d86ecc072c25502589fdbc67372166dae51aa2";
type REG is array(0 to 3) of STD_LOGIC_VECTOR (15 downto 0);
type RAMTYPE is array(0 to 8*1024-1) of STD_LOGIC_VECTOR (15 downto 0);
-- Programmspeicher 0000H-1FFFH
signal ProgRAM: RAMTYPE:=(

  x"4010",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 0000-000F
  x"4760",x"A003",x"447D",x"A003",x"4000",x"A003",x"4000",x"A003",x"4000",x"A003",x"4000",x"A003",x"4000",x"A003",x"0010",x"A003", -- 0010-001F
  x"0000",x"3000",x"0001",x"4773",x"0029",x"45E4",x"B200",x"A003",x"FFF8",x"3002",x"0001",x"4773",x"0000",x"2F10",x"A009",x"A003", -- 0020-002F
  x"FFF8",x"3004",x"0001",x"4781",x"0001",x"2F10",x"A009",x"A003",x"FFF8",x"3006",x"0007",x"4773",x"0020",x"45E4",x"465E",x"469E", -- 0030-003F
  x"B300",x"46A7",x"A003",x"FFF5",x"300E",x"0004",x"4781",x"B412",x"1000",x"A002",x"B412",x"B300",x"A003",x"FFF6",x"3013",x"0003", -- 0040-004F
  x"4781",x"B501",x"A00F",x"9001",x"A000",x"A003",x"FFF7",x"3017",x"0004",x"4781",x"B501",x"4051",x"0004",x"0000",x"4047",x"A008", -- 0050-005F
  x"9002",x"0111",x"43C2",x"4300",x"A003",x"FFF1",x"301C",x"000B",x"477A",x"42CF",x"A00A",x"2F10",x"A00A",x"9001",x"405A",x"A003", -- 0060-006F
  x"FFF5",x"3028",x"0008",x"4781",x"46B1",x"4068",x"4300",x"476B",x"A003",x"FFF7",x"3031",x"0006",x"4069",x"2800",x"FFFB",x"3038", -- 0070-007F
  x"0002",x"4069",x"2801",x"FFFB",x"303B",x"0002",x"4069",x"2802",x"FFFB",x"303E",x"0002",x"4069",x"2803",x"FFFB",x"3041",x"0004", -- 0080-008F
  x"4069",x"2F00",x"FFFB",x"3046",x"0009",x"4069",x"2F01",x"FFFB",x"3050",x"0003",x"4069",x"2F02",x"FFFB",x"3054",x"0007",x"4069", -- 0090-009F
  x"2F03",x"FFFB",x"305C",x"0007",x"4069",x"2F04",x"FFFB",x"3064",x"0004",x"4069",x"2F05",x"FFFB",x"3069",x"0007",x"4069",x"2F06", -- 00A0-00AF
  x"FFFB",x"3071",x"0004",x"4069",x"2F07",x"FFFB",x"3076",x"0004",x"4069",x"2F08",x"FFFB",x"307B",x"0003",x"4069",x"2F09",x"FFFB", -- 00B0-00BF
  x"307F",x"0003",x"4069",x"2F0A",x"FFFB",x"3083",x"0003",x"4069",x"2F0B",x"FFFB",x"3087",x"0003",x"4069",x"2F0C",x"FFFB",x"308B", -- 00C0-00CF
  x"0003",x"4069",x"2F0D",x"FFFB",x"308F",x"0007",x"4069",x"2F0E",x"FFFB",x"3097",x"0002",x"4069",x"2F0F",x"FFFB",x"309A",x"0004", -- 00D0-00DF
  x"4069",x"2F10",x"FFFB",x"309F",x"0003",x"4069",x"2F11",x"FFFB",x"30A3",x"0004",x"4069",x"2F12",x"FFFB",x"30A8",x"0005",x"4069", -- 00E0-00EF
  x"2F13",x"FFFB",x"30AE",x"0006",x"4069",x"2F14",x"FFFB",x"30B5",x"0003",x"4069",x"2F15",x"FFFB",x"30B9",x"0005",x"4069",x"2F16", -- 00F0-00FF
  x"FFFB",x"30BF",x"000C",x"4069",x"2F17",x"FFFB",x"30CC",x"0007",x"4069",x"01CB",x"FFFB",x"30D4",x"0006",x"4781",x"000A",x"0003", -- 0100-010F
  x"4047",x"A003",x"FFF8",x"30DB",x"0008",x"477A",x"42CF",x"2F10",x"A00A",x"9003",x"A00A",x"4300",x"8001",x"430B",x"A003",x"FFF3", -- 0110-011F
  x"30E4",x"0005",x"4781",x"46B1",x"4115",x"4300",x"410E",x"4300",x"476B",x"A003",x"FFF5",x"30EA",x"0005",x"4116",x"A000",x"A003", -- 0120-012F
  x"FFFA",x"30F0",x"0002",x"4116",x"A001",x"A003",x"FFFA",x"30F3",x"0002",x"4116",x"A002",x"A003",x"FFFA",x"30F6",x"0002",x"4116", -- 0130-013F
  x"A00D",x"A003",x"FFFA",x"30F9",x"0003",x"4116",x"A00F",x"A003",x"FFFA",x"30FD",x"0008",x"4116",x"A005",x"A003",x"FFFA",x"3106", -- 0140-014F
  x"0003",x"4116",x"A00B",x"A003",x"FFFA",x"310A",x"0003",x"4116",x"A008",x"A003",x"FFFA",x"310E",x"0002",x"4116",x"A00E",x"A003", -- 0150-015F
  x"FFFA",x"3111",x"0002",x"4116",x"A007",x"A003",x"FFFA",x"3114",x"0001",x"4116",x"A009",x"A003",x"FFFA",x"3116",x"0001",x"4116", -- 0160-016F
  x"A00A",x"A003",x"FFFA",x"3118",x"0004",x"4116",x"B412",x"A003",x"FFFA",x"311D",x"0004",x"4116",x"B502",x"A003",x"FFFA",x"3122", -- 0170-017F
  x"0003",x"4116",x"B501",x"A003",x"FFFA",x"3126",x"0003",x"4116",x"B434",x"A003",x"FFFA",x"312A",x"0004",x"4116",x"B300",x"A003", -- 0180-018F
  x"FFFA",x"312F",x"0005",x"4116",x"B43C",x"A003",x"FFFA",x"3135",x"0005",x"4116",x"B60C",x"A003",x"FFFA",x"313B",x"0004",x"4116", -- 0190-019F
  x"B603",x"A003",x"FFFA",x"3140",x"0005",x"4116",x"B200",x"A003",x"FFFA",x"3146",x"0004",x"4116",x"8000",x"A003",x"FFFA",x"314B", -- 01A0-01AF
  x"0002",x"4781",x"2F13",x"A00A",x"A009",x"0001",x"2F13",x"42C4",x"A003",x"FFF5",x"314E",x"0002",x"4781",x"2F13",x"A00A",x"405A", -- 01B0-01BF
  x"B501",x"4300",x"B412",x"B501",x"A00A",x"41B2",x"4286",x"B412",x"428D",x"B501",x"A00D",x"9FF6",x"B200",x"0020",x"41B2",x"A003", -- 01C0-01CF
  x"FFE9",x"3151",x"0007",x"477A",x"45E4",x"2F10",x"A00A",x"9003",x"41BD",x"42CF",x"46A7",x"A003",x"FFF4",x"3159",x"0005",x"4781", -- 01D0-01DF
  x"46B1",x"0001",x"2F10",x"A009",x"4300",x"41D3",x"FFFF",x"2F15",x"42C4",x"A003",x"FFF2",x"315F",x"0001",x"0022",x"41D4",x"A003", -- 01E0-01EF
  x"FFFA",x"3161",x"0002",x"0022",x"41D4",x"433C",x"A003",x"FFF9",x"3164",x"0004",x"4781",x"2F0F",x"A00A",x"A003",x"FFF9",x"3169", -- 01F0-01FF
  x"0005",x"4781",x"0008",x"A003",x"FFFA",x"316F",x"0006",x"4781",x"0009",x"A003",x"FFFA",x"3176",x"0006",x"4781",x"0000",x"1000", -- 0200-020F
  x"B434",x"A002",x"B412",x"B300",x"B412",x"0FFF",x"A008",x"A00E",x"A003",x"FFF1",x"317D",x"0005",x"4781",x"2F0F",x"42C4",x"A003", -- 0210-021F
  x"FFF9",x"3183",x"0007",x"4781",x"41FB",x"4286",x"4294",x"4202",x"420E",x"4300",x"A003",x"FFF5",x"318B",x"0008",x"4781",x"41FB", -- 0220-022F
  x"4286",x"4294",x"4208",x"420E",x"4300",x"A003",x"FFF5",x"3194",x"0005",x"4773",x"41FB",x"A003",x"FFFA",x"319A",x"0005",x"4773", -- 0230-023F
  x"4224",x"A003",x"FFFA",x"31A0",x"0005",x"4773",x"422F",x"A003",x"FFFA",x"31A6",x"0002",x"4773",x"4208",x"0001",x"421D",x"41FB", -- 0240-024F
  x"A003",x"FFF7",x"31A9",x"0006",x"4773",x"41FB",x"B502",x"4294",x"B434",x"420E",x"B412",x"428D",x"A009",x"A003",x"FFF3",x"31B0", -- 0250-025F
  x"0004",x"4773",x"0001",x"421D",x"4254",x"4202",x"41FB",x"A003",x"FFF6",x"31B5",x"0005",x"4773",x"424B",x"A003",x"FFFA",x"31BB", -- 0260-026F
  x"0006",x"4773",x"B434",x"423F",x"4254",x"A003",x"FFF8",x"31C2",x"0002",x"4781",x"A00A",x"A003",x"FFFA",x"31C5",x"0002",x"4781", -- 0270-027F
  x"A009",x"A003",x"FFFA",x"31C8",x"0002",x"4781",x"0001",x"A007",x"A003",x"FFF9",x"31CB",x"0002",x"4781",x"FFFF",x"A007",x"A003", -- 0280-028F
  x"FFF9",x"31CE",x"0002",x"4781",x"A000",x"A007",x"A003",x"FFF9",x"31D1",x"0001",x"4781",x"4294",x"A00D",x"A003",x"FFF9",x"31D3", -- 0290-029F
  x"0002",x"4781",x"4294",x"A00F",x"A003",x"FFF9",x"31D6",x"0001",x"4781",x"B412",x"42A2",x"A003",x"FFF9",x"31D8",x"0002",x"4781", -- 02A0-02AF
  x"0000",x"B434",x"B434",x"A002",x"B412",x"B300",x"A003",x"FFF5",x"31DB",x"0003",x"4781",x"31DF",x"0004",x"41F5",x"8FFC",x"A003", -- 02B0-02BF
  x"FFF7",x"31E4",x"0002",x"4781",x"B412",x"B502",x"A00A",x"A007",x"B412",x"A009",x"A003",x"FFF5",x"31E7",x"0002",x"4781",x"2802", -- 02C0-02CF
  x"A00A",x"4286",x"A00A",x"2802",x"A00A",x"4286",x"2802",x"B603",x"A00A",x"A00A",x"B412",x"A009",x"A009",x"A003",x"FFED",x"31EA", -- 02D0-02DF
  x"0002",x"4781",x"2802",x"A00A",x"B501",x"428D",x"2802",x"B603",x"A00A",x"A00A",x"B412",x"B501",x"428D",x"2802",x"A009",x"A009", -- 02E0-02EF
  x"A009",x"A009",x"A003",x"FFEB",x"31ED",x"0001",x"4781",x"2802",x"A00A",x"4286",x"A00A",x"A003",x"FFF7",x"31EF",x"0001",x"4781", -- 02F0-02FF
  x"2F0F",x"A00A",x"A009",x"0001",x"2F0F",x"42C4",x"A003",x"FFF5",x"31F1",x"0007",x"4781",x"2803",x"A009",x"A003",x"FFF9",x"31F9", -- 0300-030F
  x"0003",x"4781",x"5324",x"44AC",x"A00B",x"9002",x"B300",x"8FFA",x"A003",x"FFF5",x"31FD",x"0004",x"4781",x"014C",x"430B",x"A003", -- 0310-031F
  x"FFF9",x"3202",x"0005",x"4781",x"0000",x"B412",x"0010",x"A002",x"B412",x"A003",x"FFF6",x"3208",x"0003",x"4781",x"B501",x"000A", -- 0320-032F
  x"42A2",x"9001",x"8002",x"0007",x"A007",x"0030",x"A007",x"A003",x"FFF2",x"320C",x"0004",x"4781",x"B501",x"9008",x"B412",x"B501", -- 0330-033F
  x"427A",x"431D",x"4286",x"B412",x"428D",x"8FF6",x"B200",x"A003",x"FFF0",x"3211",x"0003",x"4781",x"4324",x"432E",x"431D",x"4324", -- 0340-034F
  x"432E",x"431D",x"4324",x"432E",x"431D",x"4324",x"432E",x"431D",x"B300",x"A003",x"FFEE",x"3215",x"0002",x"4781",x"434C",x"0020", -- 0350-035F
  x"431D",x"A003",x"FFF8",x"3218",x"0002",x"4781",x"A00A",x"435E",x"A003",x"FFF9",x"321B",x"0002",x"4781",x"2F07",x"A00A",x"2F0F", -- 0360-036F
  x"A00A",x"4294",x"2F10",x"A00A",x"A00D",x"A00B",x"A00E",x"2F00",x"A00A",x"A00D",x"A00B",x"A008",x"9028",x"003C",x"431D",x"321E", -- 0370-037F
  x"0003",x"41F5",x"2F07",x"A00A",x"435E",x"2F06",x"A00A",x"435E",x"003C",x"431D",x"3222",x"0004",x"41F5",x"003C",x"431D",x"3227", -- 0380-038F
  x"0003",x"41F5",x"2F0F",x"A00A",x"435E",x"2F13",x"A00A",x"435E",x"003C",x"431D",x"322B",x"0004",x"41F5",x"2F0F",x"A00A",x"2F07", -- 0390-039F
  x"A009",x"2F13",x"A00A",x"2F06",x"A009",x"000A",x"431D",x"A003",x"FFC1",x"3230",x"000A",x"4781",x"A003",x"FFFB",x"323B",x"0007", -- 03A0-03AF
  x"4781",x"436D",x"3243",x"0019",x"41F5",x"0020",x"431D",x"0008",x"431D",x"4312",x"001B",x"429B",x"9FF8",x"A003",x"FFEF",x"325D", -- 03B0-03BF
  x"0005",x"4781",x"5842",x"A003",x"A009",x"0000",x"2F10",x"A009",x"436D",x"2F0A",x"A00A",x"2F0C",x"A00A",x"2F0A",x"A00A",x"4294", -- 03C0-03CF
  x"428D",x"433C",x"3263",x"0003",x"41F5",x"3267",x"000A",x"41EF",x"46C6",x"436D",x"3272",x"0016",x"41F5",x"435E",x"43B1",x"4713", -- 03D0-03DF
  x"A003",x"FFDD",x"3289",x"0004",x"4781",x"2801",x"A00A",x"2F15",x"A009",x"A003",x"FFF7",x"328E",x"0004",x"4781",x"2801",x"A00A", -- 03E0-03EF
  x"2F15",x"A00A",x"4294",x"9002",x"0009",x"43C2",x"A003",x"FFF3",x"3293",x"0005",x"4781",x"4286",x"2F17",x"A00A",x"B502",x"4294", -- 03F0-03FF
  x"B501",x"2F17",x"A009",x"A009",x"A003",x"FFF2",x"3299",x"0009",x"4781",x"2F17",x"A00A",x"B501",x"A00A",x"A007",x"2F17",x"A009", -- 0400-040F
  x"A003",x"FFF4",x"32A3",x"0002",x"4781",x"2F17",x"A00A",x"4286",x"A003",x"FFF8",x"32A6",x"0002",x"4781",x"2F17",x"A00A",x"0002", -- 0410-041F
  x"A007",x"A003",x"FFF7",x"32A9",x"0002",x"4781",x"2F17",x"A00A",x"0003",x"A007",x"A003",x"FFF7",x"32AC",x"0002",x"4781",x"2F17", -- 0420-042F
  x"A00A",x"0004",x"A007",x"A003",x"FFF7",x"32AF",x"0002",x"4781",x"2F17",x"A00A",x"0005",x"A007",x"A003",x"FFF7",x"32B2",x"0002", -- 0430-043F
  x"4781",x"2F17",x"A00A",x"0006",x"A007",x"A003",x"FFF7",x"32B5",x"0002",x"4781",x"2F17",x"A00A",x"0007",x"A007",x"A003",x"FFF7", -- 0440-044F
  x"32B8",x"0002",x"4781",x"2F17",x"A00A",x"0008",x"A007",x"A003",x"FFF7",x"32BB",x"0001",x"4773",x"0020",x"45E4",x"465E",x"469E", -- 0450-045F
  x"B300",x"4286",x"2F10",x"A00A",x"9001",x"405A",x"A003",x"FFF1",x"32BD",x"0005",x"4781",x"B501",x"A00A",x"4286",x"B501",x"03FF", -- 0460-046F
  x"A008",x"0000",x"429B",x"9002",x"FC00",x"A007",x"B412",x"A009",x"A003",x"FFEE",x"32C3",x"0007",x"4781",x"2800",x"A00A",x"B501", -- 0470-047F
  x"0008",x"42A2",x"9009",x"0018",x"A007",x"A00A",x"B501",x"9002",x"B501",x"430B",x"B300",x"8018",x"2F03",x"A00A",x"A009",x"2F03", -- 0480-048F
  x"446B",x"2F03",x"A00A",x"2F04",x"A00A",x"4294",x"03FF",x"A008",x"0080",x"42A9",x"9009",x"2F05",x"A00A",x"A00D",x"9005",x"FFFF", -- 0490-049F
  x"2F05",x"A009",x"0013",x"431D",x"0000",x"2800",x"A009",x"A003",x"FFD1",x"32CB",x"0008",x"4781",x"2F04",x"A00A",x"2F03",x"A00A", -- 04A0-04AF
  x"429B",x"9003",x"0000",x"0000",x"8018",x"2F04",x"A00A",x"A00A",x"FFFF",x"2F04",x"446B",x"2F03",x"A00A",x"2F04",x"A00A",x"4294", -- 04B0-04BF
  x"03FF",x"A008",x"0020",x"42A2",x"9008",x"2F05",x"A00A",x"9005",x"0000",x"2F05",x"A009",x"0011",x"431D",x"A003",x"FFDA",x"32D4", -- 04C0-04CF
  x"0006",x"4781",x"0005",x"43FB",x"4426",x"A009",x"441D",x"A009",x"441D",x"A00A",x"4438",x"A009",x"4312",x"B501",x"0014",x"429B", -- 04D0-04DF
  x"9004",x"B300",x"441D",x"A00A",x"427A",x"B501",x"007F",x"429B",x"9002",x"B300",x"0008",x"B501",x"0008",x"429B",x"9012",x"4438", -- 04E0-04EF
  x"A00A",x"441D",x"A00A",x"42A2",x"900C",x"FFFF",x"441D",x"42C4",x"0001",x"4426",x"42C4",x"0008",x"431D",x"0020",x"431D",x"0008", -- 04F0-04FF
  x"431D",x"B501",x"0020",x"42A2",x"9001",x"8012",x"FFFF",x"4426",x"42C4",x"4426",x"A00A",x"A00F",x"9002",x"0006",x"43C2",x"B501", -- 0500-050F
  x"431D",x"B501",x"441D",x"A00A",x"4280",x"0001",x"441D",x"42C4",x"B501",x"0020",x"42A2",x"B502",x"0008",x"429B",x"A00B",x"A008", -- 0510-051F
  x"B412",x"001B",x"429B",x"A00B",x"A008",x"4426",x"A00A",x"A00D",x"A00E",x"9FB2",x"0020",x"431D",x"4438",x"A00A",x"441D",x"A00A", -- 0520-052F
  x"4438",x"A00A",x"4294",x"B603",x"A007",x"0000",x"B412",x"4280",x"4409",x"A003",x"FF94",x"32DB",x"0005",x"4781",x"B501",x"0030", -- 0530-053F
  x"42A2",x"A00B",x"B502",x"003A",x"42A2",x"A008",x"B502",x"0041",x"42A2",x"A00B",x"A00E",x"B501",x"9015",x"B412",x"0030",x"4294", -- 0540-054F
  x"B501",x"000A",x"42A2",x"A00B",x"9002",x"0007",x"4294",x"B501",x"2F08",x"A00A",x"42A2",x"A00B",x"9004",x"B300",x"B300",x"0000", -- 0550-055F
  x"0000",x"B412",x"A003",x"FFD7",x"32E1",x"0006",x"4781",x"4E3C",x"A003",x"441D",x"A009",x"4415",x"A009",x"0000",x"441D",x"A00A", -- 0560-056F
  x"9063",x"B501",x"4426",x"A009",x"0001",x"4441",x"A009",x"FFFF",x"444A",x"A009",x"4415",x"A00A",x"4426",x"A00A",x"A007",x"427A", -- 0570-057F
  x"002B",x"429B",x"9009",x"4426",x"A00A",x"4286",x"4426",x"A009",x"0000",x"444A",x"A009",x"8016",x"4415",x"A00A",x"4426",x"A00A", -- 0580-058F
  x"A007",x"427A",x"002D",x"429B",x"900D",x"4426",x"A00A",x"4286",x"4426",x"A009",x"0000",x"444A",x"A009",x"4441",x"A00A",x"A000", -- 0590-059F
  x"4441",x"A009",x"444A",x"A00A",x"9FD2",x"4426",x"A00A",x"441D",x"A00A",x"42A2",x"9029",x"4415",x"A00A",x"4426",x"A00A",x"A007", -- 05A0-05AF
  x"427A",x"B501",x"9015",x"453E",x"A00B",x"9007",x"B300",x"441D",x"A00A",x"A000",x"441D",x"A009",x"800A",x"B412",x"2F08",x"A00A", -- 05B0-05BF
  x"42B0",x"A007",x"4426",x"A00A",x"4286",x"4426",x"A009",x"8005",x"B300",x"4426",x"A00A",x"441D",x"A009",x"4426",x"A00A",x"441D", -- 05C0-05CF
  x"A00A",x"42A2",x"A00B",x"9FD7",x"4441",x"A00A",x"A00F",x"9001",x"A000",x"4426",x"A00A",x"441D",x"A00A",x"4294",x"4409",x"A003", -- 05D0-05DF
  x"FF83",x"32E8",x"0004",x"4781",x"42E2",x"2F0C",x"A00A",x"2F0B",x"A009",x"2F0C",x"A00A",x"427A",x"42F7",x"429B",x"2F0C",x"A00A", -- 05E0-05EF
  x"2F0D",x"A00A",x"42A2",x"A008",x"9004",x"0001",x"2F0C",x"42C4",x"8FF0",x"2F0C",x"A00A",x"2F0B",x"A009",x"2F0C",x"A00A",x"427A", -- 05F0-05FF
  x"003C",x"429B",x"9004",x"2F0C",x"A00A",x"2F0D",x"A009",x"2F0C",x"A00A",x"427A",x"42F7",x"429B",x"A00B",x"2F0C",x"A00A",x"2F0D", -- 0600-060F
  x"A00A",x"42A2",x"A008",x"9004",x"0001",x"2F0C",x"42C4",x"8FE5",x"2F0B",x"A00A",x"2F0C",x"A00A",x"B502",x"4294",x"B501",x"9003", -- 0610-061F
  x"0001",x"2F0C",x"42C4",x"42CF",x"B300",x"A003",x"FFBA",x"32ED",x"0002",x"4781",x"42E2",x"B502",x"42F7",x"4294",x"9007",x"42CF", -- 0620-062F
  x"B300",x"B300",x"B300",x"B300",x"0000",x"8023",x"42CF",x"B300",x"B412",x"0000",x"B603",x"4294",x"9016",x"42E2",x"42E2",x"B502", -- 0630-063F
  x"427A",x"B502",x"427A",x"4294",x"9004",x"B300",x"B300",x"0000",x"0000",x"B501",x"9004",x"4286",x"B412",x"4286",x"B412",x"42CF", -- 0640-064F
  x"42CF",x"4286",x"8FE7",x"B200",x"B300",x"9002",x"FFFF",x"8001",x"0000",x"A003",x"FFCC",x"32F0",x"0004",x"4781",x"42E2",x"42E2", -- 0650-065F
  x"0000",x"2F11",x"A00A",x"2F01",x"A00A",x"9003",x"B501",x"A00A",x"A007",x"B501",x"4286",x"B501",x"A00A",x"B412",x"4286",x"A00A", -- 0660-066F
  x"42CF",x"42CF",x"B603",x"42E2",x"42E2",x"462A",x"9003",x"B412",x"A00D",x"B412",x"B502",x"A00D",x"B502",x"A00A",x"A00D",x"A00B", -- 0670-067F
  x"A008",x"B502",x"B501",x"A00A",x"A007",x"2F11",x"A00A",x"429B",x"A00B",x"A008",x"9004",x"B501",x"A00A",x"A007",x"8FDA",x"42CF", -- 0680-068F
  x"B300",x"42CF",x"B434",x"A00D",x"9004",x"B300",x"B300",x"0000",x"0000",x"A003",x"FFC0",x"32F5",x"0004",x"4781",x"B412",x"0003", -- 0690-069F
  x"A007",x"B412",x"A003",x"FFF7",x"32FA",x"0008",x"4781",x"0004",x"0000",x"4047",x"A00E",x"4300",x"A003",x"FFF6",x"3303",x"0006", -- 06A0-06AF
  x"4781",x"43E5",x"2F0F",x"A00A",x"2F11",x"A00A",x"B502",x"4294",x"4300",x"2F11",x"A009",x"0020",x"45E4",x"41BD",x"0001",x"2F01", -- 06B0-06BF
  x"A009",x"A003",x"FFEB",x"330A",x"0009",x"4781",x"2F0A",x"A00A",x"42E2",x"2F0B",x"A00A",x"42E2",x"2F0C",x"A00A",x"42E2",x"2F0D", -- 06C0-06CF
  x"A00A",x"42E2",x"B502",x"A007",x"2F0D",x"A009",x"B501",x"2F0A",x"A009",x"B501",x"2F0B",x"A009",x"2F0C",x"A009",x"0020",x"45E4", -- 06D0-06DF
  x"B501",x"901F",x"B603",x"465E",x"B501",x"9009",x"42E2",x"42E2",x"B200",x"42CF",x"42CF",x"469E",x"B300",x"430B",x"8011",x"B200", -- 06E0-06EF
  x"B603",x"4567",x"9005",x"B200",x"B300",x"0003",x"43C2",x"8008",x"B434",x"B300",x"B412",x"B300",x"2F10",x"A00A",x"9001",x"405A", -- 06F0-06FF
  x"8FDD",x"B200",x"42CF",x"2F0D",x"A009",x"42CF",x"2F0C",x"A009",x"42CF",x"2F0B",x"A009",x"42CF",x"2F0A",x"A009",x"A003",x"FFB3", -- 0700-070F
  x"3314",x"0004",x"4781",x"2F02",x"A00A",x"2802",x"A009",x"2F00",x"A00A",x"9006",x"003C",x"431D",x"3319",x"0004",x"41F5",x"8003", -- 0710-071F
  x"331E",x"0002",x"41F5",x"436D",x"2F09",x"A00A",x"0100",x"44D2",x"B502",x"A00A",x"003C",x"429B",x"9002",x"B200",x"802B",x"2F00", -- 0720-072F
  x"A00A",x"900C",x"003C",x"431D",x"3321",x"0003",x"41F5",x"46C6",x"003C",x"431D",x"3325",x"0004",x"41F5",x"801C",x"001B",x"431D", -- 0730-073F
  x"005B",x"431D",x"0033",x"431D",x"0036",x"431D",x"006D",x"431D",x"46C6",x"2F10",x"A00A",x"A00D",x"9003",x"332A",x"0002",x"41F5", -- 0740-074F
  x"001B",x"431D",x"005B",x"431D",x"0033",x"431D",x"0039",x"431D",x"006D",x"431D",x"8FC8",x"A003",x"FFB3",x"332D",x"0005",x"4781", -- 0750-075F
  x"3333",x"000B",x"41F5",x"436D",x"436D",x"4713",x"A003",x"FFF5",x"333F",x"0006",x"4781",x"0000",x"2F01",x"A009",x"A003",x"FFF8", -- 0760-076F
  x"3346",x"000C",x"4781",x"42CF",x"42E2",x"A003",x"FFF9",x"3353",x"000A",x"4781",x"42CF",x"46A7",x"A003",x"FFF9",x"335E",x"0003", -- 0770-077F
  x"4781",x"42CF",x"2F10",x"A00A",x"9002",x"46A7",x"8001",x"42E2",x"A003",x"FFF4",x"3362",x"000A",x"4781",x"46B1",x"0001",x"2F10", -- 0780-078F
  x"A009",x"4772",x"A003",x"FFF6",x"336D",x"0008",x"4781",x"46B1",x"0001",x"2F10",x"A009",x"4779",x"A003",x"FFF6",x"3376",x"0001", -- 0790-079F
  x"4781",x"46B1",x"0001",x"2F10",x"A009",x"4780",x"A003",x"FFF6",x"3378",x"0001",x"4773",x"0000",x"2F10",x"A009",x"43EE",x"410E", -- 07A0-07AF
  x"4300",x"476B",x"A003",x"FFF4",x"337A",x"0003",x"4781",x"2F16",x"A00A",x"9005",x"4324",x"B300",x"4324",x"B300",x"8006",x"4324", -- 07B0-07BF
  x"432E",x"431D",x"4324",x"432E",x"431D",x"4324",x"432E",x"431D",x"4324",x"432E",x"431D",x"B300",x"A003",x"FFE6",x"337E",x"0003", -- 07C0-07CF
  x"4781",x"3382",x"0001",x"41F5",x"0022",x"431D",x"47B7",x"0022",x"431D",x"3384",x"0001",x"41F5",x"A003",x"FFF0",x"3386",x"0005", -- 07D0-07DF
  x"4781",x"2F16",x"A009",x"2F00",x"A00A",x"42E2",x"0000",x"2F00",x"A009",x"338C",x"0008",x"41EF",x"46C6",x"0004",x"0000",x"4047", -- 07E0-07EF
  x"A00E",x"0010",x"A009",x"436D",x"003C",x"431D",x"3395",x"0006",x"41F5",x"436D",x"339C",x"0002",x"41F5",x"0000",x"B603",x"A007", -- 07F0-07FF
  x"B501",x"2F03",x"429B",x"9002",x"B300",x"2F04",x"B501",x"2F17",x"429B",x"9005",x"B300",x"2D00",x"2F80",x"A009",x"2F80",x"B501", -- 0800-080F
  x"2F05",x"429B",x"9002",x"B300",x"2F00",x"A00A",x"47D1",x"4286",x"B501",x"0010",x"429B",x"9FE2",x"B300",x"339F",x"0004",x"41F5", -- 0810-081F
  x"B501",x"434C",x"33A4",x"0001",x"41F5",x"B501",x"000F",x"A007",x"434C",x"0010",x"A007",x"B603",x"42A9",x"A00B",x"9FCA",x"B200", -- 0820-082F
  x"436D",x"003C",x"431D",x"33A6",x"0007",x"41F5",x"42CF",x"2F00",x"A009",x"A003",x"FFA3",x"33AE",x"0005",x"4069",x"2F20",x"FFFB", -- 0830-083F
  x"33B4",x"0008",x"4781",x"2F20",x"A00A",x"B501",x"4074",x"B501",x"4286",x"2F20",x"A009",x"A009",x"A003",x"FFF2",x"33BD",x"0004", -- 0840-084F
  x"4781",x"B501",x"900D",x"B434",x"B434",x"B502",x"A00A",x"B502",x"A009",x"B412",x"4286",x"B412",x"4286",x"B434",x"428D",x"8FF1", -- 0850-085F
  x"B300",x"B200",x"A003",x"FFEA",x"33C2",x"0004",x"4781",x"B434",x"B434",x"B501",x"9008",x"B434",x"B434",x"B603",x"A009",x"4286", -- 0860-086F
  x"B434",x"428D",x"8FF6",x"B300",x"B200",x"A003",x"FFED",x"33C7",x"0004",x"4781",x"B412",x"B501",x"A00A",x"435E",x"4286",x"B412", -- 0870-087F
  x"428D",x"B501",x"A00D",x"9FF6",x"B200",x"A003",x"FFF0",x"33CC",x"0003",x"4781",x"B603",x"42A2",x"9001",x"B412",x"B300",x"A003", -- 0880-088F
  x"FFF6",x"33D0",x"0003",x"4781",x"B603",x"42A9",x"9001",x"B412",x"B300",x"A003",x"FFF6",x"33D4",x"0006",x"4116",x"A017",x"A003", -- 0890-089F
  x"FFFA",x"33DB",x"0007",x"4116",x"A018",x"A003",x"FFFA",x"33E3",x"0009",x"4781",x"42E2",x"A017",x"A018",x"9FFD",x"42CF",x"B300", -- 08A0-08AF
  x"A003",x"FFF5",x"33ED",x"0001",x"4069",x"1401",x"FFFB",x"33EF",x"0001",x"4069",x"1601",x"FFFB",x"33F1",x"0001",x"4069",x"1801", -- 08B0-08BF
  x"FFFB",x"33F3",x"0004",x"4781",x"0007",x"43FB",x"444A",x"A009",x"4441",x"A009",x"4438",x"A009",x"442F",x"A009",x"4426",x"A009", -- 08C0-08CF
  x"441D",x"A009",x"4415",x"A009",x"4415",x"A00A",x"442F",x"A00A",x"9001",x"A00B",x"441D",x"A00A",x"4438",x"A00A",x"A007",x"4286", -- 08D0-08DF
  x"444A",x"A00A",x"B502",x"0000",x"4867",x"444A",x"A00A",x"B501",x"4426",x"A00A",x"441D",x"A00A",x"0000",x"B60C",x"A00A",x"B434", -- 08E0-08EF
  x"B434",x"4441",x"A00A",x"4438",x"A00A",x"48AA",x"B300",x"A009",x"B300",x"B434",x"4286",x"B434",x"4286",x"B434",x"428D",x"B501", -- 08F0-08FF
  x"A00D",x"9FEA",x"B300",x"B200",x"4409",x"A003",x"FFBA",x"33F8",x"0006",x"4781",x"0007",x"43FB",x"444A",x"A009",x"4441",x"A009", -- 0900-090F
  x"4438",x"A009",x"442F",x"A009",x"4426",x"A009",x"441D",x"A009",x"4415",x"A009",x"4415",x"A00A",x"441D",x"A00A",x"4438",x"A00A", -- 0910-091F
  x"488A",x"4286",x"444A",x"A00A",x"4415",x"A00A",x"442F",x"A00A",x"429B",x"903B",x"0000",x"441D",x"A00A",x"4438",x"A00A",x"488A", -- 0920-092F
  x"0000",x"B434",x"B502",x"B501",x"441D",x"A00A",x"42A2",x"9009",x"4426",x"A00A",x"B501",x"A00A",x"B412",x"4286",x"4426",x"A009", -- 0930-093F
  x"8001",x"0000",x"B412",x"4438",x"A00A",x"42A2",x"9009",x"4441",x"A00A",x"B501",x"A00A",x"B412",x"4286",x"4441",x"A009",x"8001", -- 0940-094F
  x"0000",x"A001",x"444A",x"A00A",x"B501",x"4286",x"444A",x"A009",x"A009",x"B434",x"B434",x"4286",x"B603",x"4294",x"A00D",x"9FD1", -- 0950-095F
  x"B200",x"444A",x"A00A",x"A009",x"8063",x"B412",x"0001",x"4294",x"B412",x"0001",x"441D",x"A00A",x"4438",x"A00A",x"488A",x"0000", -- 0960-096F
  x"B434",x"B502",x"B501",x"441D",x"A00A",x"42A2",x"9009",x"4426",x"A00A",x"B501",x"A00A",x"B412",x"4286",x"4426",x"A009",x"8001", -- 0970-097F
  x"0000",x"B412",x"4438",x"A00A",x"42A2",x"900A",x"4441",x"A00A",x"B501",x"A00A",x"B412",x"4286",x"4441",x"A009",x"A00B",x"8001", -- 0980-098F
  x"FFFF",x"A001",x"444A",x"A00A",x"B501",x"4286",x"444A",x"A009",x"A009",x"B434",x"B434",x"4286",x"B603",x"4294",x"A00D",x"9FD0", -- 0990-099F
  x"B200",x"A00D",x"9025",x"B501",x"444A",x"A009",x"B434",x"A00B",x"B434",x"B434",x"0001",x"441D",x"A00A",x"4438",x"A00A",x"488A", -- 09A0-09AF
  x"0000",x"B434",x"0000",x"444A",x"A00A",x"A00A",x"A00B",x"A001",x"444A",x"A00A",x"B501",x"4286",x"444A",x"A009",x"A009",x"B434", -- 09B0-09BF
  x"B434",x"4286",x"B603",x"4294",x"A00D",x"9FEB",x"B200",x"B300",x"4409",x"A003",x"FF3C",x"33FF",x"0004",x"4116",x"A014",x"A003", -- 09C0-09CF
  x"FFFA",x"3404",x"0005",x"4781",x"0010",x"42E2",x"A014",x"42CF",x"428D",x"B501",x"A00D",x"9FF9",x"B200",x"A003",x"FFF2",x"340A", -- 09D0-09DF
  x"0005",x"4781",x"0000",x"B434",x"B434",x"49D4",x"A003",x"FFF7",x"3410",x"0004",x"4781",x"0007",x"43FB",x"444A",x"A009",x"4441", -- 09E0-09EF
  x"A009",x"4438",x"A009",x"442F",x"A009",x"4426",x"A009",x"441D",x"A009",x"4415",x"A009",x"441D",x"A00A",x"4438",x"A00A",x"42A2", -- 09F0-09FF
  x"900A",x"4415",x"A00A",x"441D",x"A00A",x"4426",x"A00A",x"0000",x"0000",x"0000",x"80D9",x"441D",x"A00A",x"0000",x"4426",x"A00A", -- 0A00-0A0F
  x"B502",x"A007",x"A00A",x"A00B",x"B502",x"444A",x"A00A",x"A007",x"A009",x"4286",x"B603",x"4294",x"A00D",x"9FF0",x"B200",x"444A", -- 0A10-0A1F
  x"A00A",x"441D",x"A00A",x"A007",x"4438",x"A00A",x"4294",x"4426",x"A009",x"FFFF",x"444A",x"A00A",x"441D",x"A00A",x"A007",x"A009", -- 0A20-0A2F
  x"0001",x"441D",x"42C4",x"441D",x"A00A",x"4438",x"A00A",x"4294",x"0000",x"4426",x"A00A",x"4438",x"A00A",x"A007",x"A00A",x"A00B", -- 0A30-0A3F
  x"4426",x"A00A",x"4438",x"A00A",x"A007",x"428D",x"A00A",x"A00B",x"4441",x"A00A",x"4438",x"A00A",x"A007",x"428D",x"A00A",x"49D4", -- 0A40-0A4F
  x"B412",x"B300",x"B501",x"4426",x"A00A",x"4438",x"A00A",x"A007",x"4286",x"A009",x"0000",x"4426",x"A00A",x"4441",x"A00A",x"4438", -- 0A50-0A5F
  x"A00A",x"48AA",x"B200",x"B412",x"B300",x"0000",x"4426",x"A00A",x"4438",x"A00A",x"A007",x"A00A",x"A001",x"4426",x"A00A",x"4438", -- 0A60-0A6F
  x"A00A",x"A007",x"A009",x"902B",x"0001",x"4438",x"A00A",x"0000",x"B434",x"B502",x"4426",x"A00A",x"B502",x"A007",x"A00A",x"B412", -- 0A70-0A7F
  x"4441",x"A00A",x"A007",x"A00A",x"A00B",x"A001",x"B412",x"42E2",x"B502",x"4426",x"A00A",x"A007",x"A009",x"42CF",x"B434",x"B434", -- 0A80-0A8F
  x"4286",x"B603",x"4294",x"A00D",x"9FE3",x"B200",x"FFFF",x"4426",x"A00A",x"4438",x"A00A",x"A007",x"4286",x"42C4",x"8FD4",x"FFFF", -- 0A90-0A9F
  x"4426",x"42C4",x"4286",x"B603",x"4294",x"A00D",x"9F92",x"B200",x"4438",x"A00A",x"0000",x"444A",x"A00A",x"B502",x"A007",x"A00A", -- 0AA0-0AAF
  x"A00B",x"B502",x"444A",x"A00A",x"A007",x"A009",x"4286",x"B603",x"4294",x"A00D",x"9FF0",x"B200",x"4438",x"A00A",x"444A",x"A00A", -- 0AB0-0ABF
  x"428D",x"A009",x"441D",x"A00A",x"4438",x"A00A",x"4294",x"444A",x"A00A",x"4438",x"A00A",x"A007",x"A009",x"4415",x"A00A",x"4438", -- 0AC0-0ACF
  x"A00A",x"444A",x"A00A",x"4415",x"A00A",x"442F",x"A00A",x"9001",x"A00B",x"441D",x"A00A",x"4438",x"A00A",x"4294",x"444A",x"A00A", -- 0AD0-0ADF
  x"4438",x"A00A",x"A007",x"4286",x"4409",x"A003",x"FF01",x"3415",x"0008",x"4069",x"2F21",x"FFFB",x"341E",x"0008",x"4069",x"2F22", -- 0AE0-0AEF
  x"FFFB",x"3427",x"0008",x"4069",x"2F23",x"FFFB",x"3430",x"000E",x"4069",x"2F24",x"FFFB",x"343F",x"000C",x"4069",x"2F25",x"FFFB", -- 0AF0-0AFF
  x"344C",x"0006",x"4069",x"2F26",x"FFFB",x"3453",x"0004",x"4069",x"2F27",x"FFFB",x"3458",x"0004",x"4781",x"B412",x"B603",x"A007", -- 0B00-0B0F
  x"428D",x"B502",x"A00D",x"A00B",x"B502",x"A00A",x"A00D",x"A008",x"9005",x"B412",x"428D",x"B412",x"428D",x"8FF3",x"B300",x"B412", -- 0B10-0B1F
  x"A003",x"FFE8",x"345D",x"0012",x"4781",x"428D",x"B412",x"B502",x"A009",x"0004",x"0000",x"4047",x"A00E",x"B412",x"9001",x"A000", -- 0B20-0B2F
  x"A003",x"FFF0",x"3470",x"000D",x"4781",x"B502",x"9015",x"B502",x"0001",x"429B",x"B502",x"A00A",x"000C",x"0000",x"4047",x"A008", -- 0B30-0B3F
  x"A00D",x"A008",x"9007",x"A00A",x"B412",x"B300",x"B412",x"9001",x"A000",x"8001",x"4B25",x"8003",x"B200",x"B300",x"0000",x"A003", -- 0B40-0B4F
  x"FFE1",x"347E",x"000C",x"4781",x"B501",x"A00A",x"B501",x"A00F",x"9003",x"A000",x"FFFF",x"8001",x"0000",x"B434",x"B434",x"B501", -- 0B50-0B5F
  x"0004",x"0000",x"4047",x"A008",x"900E",x"B412",x"B300",x"2F27",x"A00A",x"9002",x"FFFF",x"8001",x"3FFF",x"A008",x"B501",x"A00A", -- 0B60-0B6F
  x"B412",x"4286",x"8004",x"B502",x"A009",x"0001",x"B412",x"A003",x"FFD8",x"348B",x"000D",x"4781",x"B501",x"2F25",x"A00A",x"42A2", -- 0B70-0B7F
  x"A00B",x"9006",x"3499",x"0004",x"41EF",x"46C6",x"0369",x"43C2",x"2F23",x"A009",x"A003",x"FFED",x"349E",x"000B",x"4781",x"2F23", -- 0B80-0B8F
  x"A00A",x"B603",x"A009",x"4286",x"B603",x"A007",x"4B7C",x"B603",x"B412",x"0000",x"4867",x"B412",x"B300",x"A003",x"FFED",x"34AA", -- 0B90-0B9F
  x"0010",x"4781",x"2F22",x"A009",x"2F21",x"A009",x"2F21",x"4B54",x"B502",x"42E2",x"2F22",x"4B54",x"B502",x"42CF",x"A007",x"4286", -- 0BA0-0BAF
  x"4B8F",x"A003",x"FFEC",x"34BB",x"0001",x"4781",x"4BA2",x"490A",x"4B0D",x"4B35",x"A003",x"FFF7",x"34BD",x"0001",x"4781",x"A000", -- 0BB0-0BBF
  x"4BB6",x"A003",x"FFF9",x"34BF",x"0001",x"4781",x"4BA2",x"48C4",x"4B0D",x"4B35",x"A003",x"FFF7",x"34C1",x"0007",x"4773",x"2F11", -- 0BC0-0BCF
  x"A00A",x"0004",x"A007",x"46A7",x"A003",x"FFF6",x"34C9",x"0004",x"4781",x"B501",x"A00D",x"9002",x"0000",x"43C2",x"B501",x"2F21", -- 0BD0-0BDF
  x"A009",x"2F21",x"4B54",x"B434",x"B300",x"B502",x"A007",x"428D",x"A00A",x"B412",x"0001",x"42A9",x"9018",x"0001",x"B502",x"A00F", -- 0BE0-0BEF
  x"A00B",x"9007",x"B412",x"B501",x"A007",x"B412",x"B501",x"4BB6",x"8FF5",x"B412",x"B300",x"B501",x"2F26",x"A009",x"B434",x"B502", -- 0BF0-0BFF
  x"4BC6",x"B434",x"B434",x"4BC6",x"8004",x"B300",x"0001",x"2F26",x"A009",x"4BA2",x"49EB",x"4B0D",x"4B35",x"42E2",x"4B0D",x"4B35", -- 0C00-0C0F
  x"42CF",x"2F26",x"A00A",x"428D",x"9007",x"B412",x"2F26",x"A00A",x"4BD9",x"B412",x"B300",x"B412",x"A003",x"FFB8",x"34CE",x"0004", -- 0C10-0C1F
  x"4781",x"0000",x"42E2",x"4324",x"B501",x"9007",x"432E",x"431D",x"42CF",x"B300",x"FFFF",x"42E2",x"8001",x"B300",x"4324",x"B501", -- 0C20-0C2F
  x"42F7",x"A00E",x"9007",x"432E",x"431D",x"42CF",x"B300",x"FFFF",x"42E2",x"8001",x"B300",x"4324",x"B501",x"42F7",x"A00E",x"9003", -- 0C30-0C3F
  x"432E",x"431D",x"8001",x"B300",x"4324",x"432E",x"431D",x"B300",x"42CF",x"B300",x"A003",x"FFD2",x"34D3",x"0001",x"4781",x"2F21", -- 0C40-0C4F
  x"A009",x"2F21",x"4B54",x"B434",x"9003",x"34D5",x"0001",x"41F5",x"B502",x"A007",x"428D",x"B501",x"A00A",x"4C21",x"B412",x"428D", -- 0C50-0C5F
  x"B412",x"B502",x"9008",x"428D",x"B501",x"A00A",x"434C",x"B412",x"428D",x"B412",x"8FF6",x"B300",x"B300",x"0020",x"431D",x"A003", -- 0C60-0C6F
  x"FFDB",x"34D7",x"0002",x"4781",x"B412",x"4C4F",x"4C4F",x"A003",x"FFF8",x"34DA",x"000B",x"4069",x"2F28",x"FFFB",x"34E6",x"0009", -- 0C70-0C7F
  x"4069",x"2F29",x"FFFB",x"34F0",x"000D",x"4781",x"2F23",x"A00A",x"A003",x"FFF9",x"34FE",x"000D",x"4781",x"2F23",x"A009",x"A003", -- 0C80-0C8F
  x"FFF9",x"350C",x"000B",x"4781",x"2F29",x"A00A",x"2F28",x"A009",x"2F23",x"A00A",x"2F29",x"A009",x"A003",x"FFF3",x"3518",x"000A", -- 0C90-0C9F
  x"4781",x"0000",x"B502",x"A009",x"B501",x"A00A",x"B412",x"FFFF",x"B502",x"A009",x"8000",x"A00A",x"4286",x"A00E",x"A00D",x"A003", -- 0CA0-0CAF
  x"FFED",x"3523",x"0004",x"4781",x"0000",x"1C00",x"0007",x"0000",x"4047",x"4CA1",x"9005",x"B200",x"FFFF",x"0007",x"0000",x"4047", -- 0CB0-0CBF
  x"0006",x"0000",x"4047",x"4CA1",x"9005",x"B200",x"FFFF",x"0006",x"0000",x"4047",x"0004",x"0000",x"4047",x"4CA1",x"9005",x"B200", -- 0CC0-0CCF
  x"FFFF",x"0004",x"0000",x"4047",x"2000",x"0005",x"0FFF",x"4047",x"4CA1",x"9004",x"B300",x"0006",x"0000",x"4047",x"0006",x"0FFF", -- 0CD0-0CDF
  x"4047",x"4CA1",x"9004",x"B300",x"0007",x"0000",x"4047",x"0007",x"07FF",x"4047",x"4CA1",x"9004",x"B300",x"0007",x"0800",x"4047", -- 0CE0-0CEF
  x"2F25",x"A009",x"2F24",x"A009",x"2F27",x"A009",x"2F24",x"A00A",x"2F23",x"A009",x"4C94",x"4C94",x"A003",x"FFB3",x"3528",x"0003", -- 0CF0-0CFF
  x"4781",x"B501",x"2F21",x"A009",x"2F21",x"4B54",x"B501",x"2F21",x"4294",x"900E",x"2F23",x"A00A",x"4286",x"B412",x"B502",x"B60C", -- 0D00-0D0F
  x"B502",x"A007",x"4B7C",x"4851",x"4B25",x"B412",x"B300",x"8002",x"B200",x"B300",x"A003",x"FFE2",x"352C",x"0003",x"4781",x"B412", -- 0D10-0D1F
  x"4D01",x"B412",x"4D01",x"A003",x"FFF7",x"3530",x"0001",x"4781",x"4C86",x"B434",x"B434",x"4BB6",x"B412",x"4C8D",x"4D01",x"A003", -- 0D20-0D2F
  x"FFF4",x"3532",x"0001",x"4781",x"4C86",x"B434",x"B434",x"4BBF",x"B412",x"4C8D",x"4D01",x"A003",x"FFF4",x"3534",x"0001",x"4781", -- 0D30-0D3F
  x"4C86",x"B434",x"B434",x"4BC6",x"B412",x"4C8D",x"4D01",x"A003",x"FFF4",x"3536",x"0001",x"4781",x"4C86",x"B434",x"B434",x"4BD9", -- 0D40-0D4F
  x"B412",x"B300",x"B412",x"4C8D",x"4D01",x"A003",x"FFF2",x"3538",x"0003",x"4781",x"4C86",x"B434",x"B434",x"4BD9",x"B300",x"B412", -- 0D50-0D5F
  x"4C8D",x"4D01",x"A003",x"FFF3",x"353C",x"0003",x"4781",x"4C86",x"B434",x"B434",x"B501",x"9004",x"B412",x"B502",x"4D5A",x"8FFA", -- 0D60-0D6F
  x"B300",x"B412",x"4C8D",x"4D01",x"A003",x"FFEE",x"3540",x"0002",x"4781",x"4C86",x"B434",x"B434",x"B603",x"4D67",x"B434",x"B502", -- 0D70-0D7F
  x"4D4C",x"B434",x"B434",x"4D4C",x"B434",x"4C8D",x"4D1F",x"A003",x"FFED",x"3543",x"0007",x"4781",x"4C86",x"B434",x"B434",x"0007", -- 0D80-0D8F
  x"43FB",x"441D",x"A009",x"4415",x"A009",x"0000",x"441D",x"A00A",x"9063",x"B501",x"4426",x"A009",x"0001",x"4441",x"A009",x"FFFF", -- 0D90-0D9F
  x"444A",x"A009",x"4415",x"A00A",x"4426",x"A00A",x"A007",x"427A",x"002B",x"429B",x"9009",x"4426",x"A00A",x"4286",x"4426",x"A009", -- 0DA0-0DAF
  x"0000",x"444A",x"A009",x"8016",x"4415",x"A00A",x"4426",x"A00A",x"A007",x"427A",x"002D",x"429B",x"900D",x"4426",x"A00A",x"4286", -- 0DB0-0DBF
  x"4426",x"A009",x"0000",x"444A",x"A009",x"4441",x"A00A",x"A000",x"4441",x"A009",x"444A",x"A00A",x"9FD2",x"4426",x"A00A",x"441D", -- 0DC0-0DCF
  x"A00A",x"42A2",x"9029",x"4415",x"A00A",x"4426",x"A00A",x"A007",x"427A",x"B501",x"9015",x"453E",x"A00B",x"9007",x"B300",x"441D", -- 0DD0-0DDF
  x"A00A",x"A000",x"441D",x"A009",x"800A",x"B412",x"2F08",x"A00A",x"4D40",x"4D28",x"4426",x"A00A",x"4286",x"4426",x"A009",x"8005", -- 0DE0-0DEF
  x"B300",x"4426",x"A00A",x"441D",x"A009",x"4426",x"A00A",x"441D",x"A00A",x"42A2",x"A00B",x"9FD7",x"4441",x"A00A",x"A00F",x"9001", -- 0DF0-0DFF
  x"A000",x"4426",x"A00A",x"441D",x"A00A",x"4294",x"B501",x"9006",x"B300",x"4415",x"A00A",x"4426",x"A00A",x"A007",x"4409",x"B434", -- 0E00-0E0F
  x"4C8D",x"B412",x"4D01",x"B412",x"A003",x"FF73",x"354B",x"0002",x"0022",x"41D4",x"4D8C",x"B300",x"A003",x"FFF8",x"354E",x"0008", -- 0E10-0E1F
  x"4781",x"43E5",x"0020",x"45E4",x"465E",x"B501",x"9011",x"469E",x"B300",x"4286",x"41FB",x"B412",x"2F0F",x"A009",x"B501",x"46A7", -- 0E20-0E2F
  x"410E",x"4300",x"2F0F",x"A009",x"0001",x"2F10",x"A009",x"8003",x"B200",x"0003",x"43C2",x"A003",x"4D8C",x"A003",x"FFDF",x"3557", -- 0E30-0E3F
  x"0001",x"4781",x"4C86",x"B434",x"B434",x"0004",x"43FB",x"B501",x"A00F",x"9002",x"0012",x"43C2",x"0002",x"442F",x"A009",x"4426", -- 0E40-0E4F
  x"A009",x"441D",x"A009",x"0001",x"4426",x"A00A",x"442F",x"A00A",x"49E2",x"4426",x"A009",x"9003",x"441D",x"A00A",x"4D40",x"4426", -- 0E50-0E5F
  x"A00A",x"9008",x"441D",x"A00A",x"441D",x"A00A",x"4D40",x"441D",x"A009",x"8FEA",x"4409",x"B412",x"4C8D",x"4D01",x"A003",x"FFCF", -- 0E60-0E6F
  x"3559",x"0001",x"4781",x"2F08",x"A00A",x"0010",x"429B",x"9002",x"4C4F",x"802C",x"4C86",x"B412",x"B501",x"A00F",x"9004",x"A000", -- 0E70-0E7F
  x"355B",x"0001",x"41F5",x"B501",x"A00D",x"9005",x"355D",x"0002",x"41F5",x"B300",x"801A",x"FFFF",x"B412",x"B501",x"9004",x"2F08", -- 0E80-0E8F
  x"A00A",x"4BD9",x"8FFA",x"B300",x"B501",x"A00F",x"A00B",x"900A",x"0030",x"A007",x"B501",x"0039",x"42A9",x"9002",x"0007",x"A007", -- 0E90-0E9F
  x"431D",x"8FF2",x"0020",x"431D",x"B300",x"4C8D",x"A003",x"FFC8",x"3560",x"0002",x"4781",x"B412",x"4E73",x"4E73",x"A003",x"FFF8", -- 0EA0-0EAF
  x"3563",x"0006",x"4781",x"2F27",x"A00A",x"9002",x"FFFF",x"8001",x"3FFF",x"A008",x"B501",x"4286",x"B412",x"A00A",x"A003",x"FFF0", -- 0EB0-0EBF
  x"356A",x"0004",x"4781",x"4051",x"B501",x"0004",x"0000",x"4047",x"42A2",x"9003",x"B300",x"0000",x"800B",x"4EB3",x"B412",x"B300", -- 0EC0-0ECF
  x"0004",x"0000",x"4047",x"42A2",x"9002",x"0000",x"8001",x"FFFF",x"A003",x"FFE6",x"356F",x"0001",x"4781",x"B502",x"4EC3",x"9011", -- 0ED0-0EDF
  x"B412",x"4EB3",x"3FFF",x"A008",x"B434",x"B603",x"42A9",x"9005",x"B412",x"B300",x"A007",x"A00A",x"8003",x"B200",x"B300",x"0000", -- 0EE0-0EEF
  x"8003",x"9002",x"B300",x"0000",x"A003",x"FFE4",x"3571",x"0001",x"4781",x"B603",x"4EDD",x"A003",x"FFF9",x"3573",x"0001",x"4781", -- 0EF0-0EFF
  x"B501",x"42E2",x"B434",x"B434",x"B502",x"4EC3",x"A00D",x"B502",x"A00D",x"A008",x"42CF",x"4EC3",x"A00D",x"A008",x"9002",x"B200", -- 0F00-0F0F
  x"8072",x"B502",x"4EC3",x"A00D",x"9017",x"B501",x"4286",x"4B8F",x"B434",x"B502",x"A009",x"0004",x"0000",x"4047",x"B502",x"428D", -- 0F10-0F1F
  x"42C4",x"B501",x"42E2",x"A007",x"A009",x"42CF",x"428D",x"0004",x"0000",x"4047",x"A00E",x"8057",x"B502",x"4EB3",x"3FFF",x"A008", -- 0F20-0F2F
  x"B434",x"B603",x"42A9",x"9008",x"B412",x"B300",x"B434",x"42E2",x"A007",x"A009",x"42CF",x"801F",x"B501",x"4286",x"4B8F",x"B412", -- 0F30-0F3F
  x"42E2",x"B501",x"42E2",x"B412",x"4851",x"B300",x"42CF",x"0004",x"0000",x"4047",x"B502",x"428D",x"A00A",x"A00E",x"B502",x"428D", -- 0F40-0F4F
  x"A009",x"B412",x"B502",x"42CF",x"A007",x"A009",x"428D",x"0004",x"0000",x"4047",x"A00E",x"4EB3",x"3FFF",x"A008",x"B603",x"A007", -- 0F50-0F5F
  x"428D",x"A00A",x"A00D",x"B502",x"0001",x"42A9",x"A008",x"9002",x"428D",x"8FF4",x"B502",x"A00A",x"4EC3",x"A00D",x"B502",x"0001", -- 0F60-0F6F
  x"429B",x"A008",x"9003",x"B300",x"A00A",x"800D",x"B412",x"428D",x"B412",x"0004",x"0000",x"4047",x"A00E",x"B502",x"A009",x"0004", -- 0F70-0F7F
  x"0000",x"4047",x"A00E",x"A003",x"FF78",x"3575",x"0001",x"4781",x"B501",x"4EC3",x"9016",x"3577",x"0002",x"41F5",x"4EB3",x"3FFF", -- 0F80-0F8F
  x"A008",x"B502",x"A007",x"B412",x"B603",x"42A9",x"9005",x"B501",x"A00A",x"4F88",x"4286",x"8FF8",x"B200",x"357A",x"0002",x"41F5", -- 0F90-0F9F
  x"8001",x"4E73",x"A003",x"FFE1",x"357D",x"0002",x"4781",x"B412",x"4F88",x"4F88",x"A003",x"FFF8",x"3580",x"0006",x"4069",x"2F2A", -- 0FA0-0FAF
  x"FFFB",x"3587",x"0001",x"4781",x"2F2A",x"A00A",x"2801",x"A00A",x"2F2A",x"A009",x"A003",x"FFF5",x"3589",x"0001",x"4781",x"0000", -- 0FB0-0FBF
  x"2801",x"A00A",x"428D",x"2F2A",x"A00A",x"4294",x"900A",x"2801",x"A00A",x"0002",x"4294",x"2F2A",x"A00A",x"4294",x"B434",x"4F00", -- 0FC0-0FCF
  x"8FEF",x"B412",x"2F2A",x"A009",x"A003",x"FFE6",x"358B",x"0005",x"4781",x"B501",x"4EC3",x"9019",x"B501",x"42E2",x"4EB3",x"3FFF", -- 0FD0-0FDF
  x"A008",x"B412",x"B502",x"A007",x"428D",x"B412",x"B501",x"900A",x"B412",x"B501",x"A00A",x"4FD9",x"B502",x"A009",x"428D",x"B412", -- 0FE0-0FEF
  x"428D",x"8FF4",x"B200",x"42CF",x"8001",x"4D01",x"A003",x"FFDE",x"3591",x"0007",x"4781",x"B501",x"4EC3",x"9028",x"4EB3",x"3FFF", -- 0FF0-0FFF
  x"A008",x"B501",x"9021",x"B412",x"436D",x"B502",x"435E",x"B501",x"435E",x"B501",x"A00A",x"B501",x"435E",x"B501",x"4051",x"3FFF", -- 1000-100F
  x"42A9",x"A00B",x"9005",x"FFFF",x"435E",x"FFFF",x"435E",x"8005",x"B501",x"4051",x"4EB3",x"435E",x"435E",x"B501",x"4F88",x"4FFB", -- 1010-101F
  x"4286",x"B412",x"428D",x"8FDD",x"B200",x"8001",x"B300",x"A003",x"FFCF",x"3599",x"000F",x"4781",x"B501",x"4EC3",x"9028",x"2F23", -- 1020-102F
  x"A00A",x"0004",x"0000",x"4047",x"A00E",x"B412",x"4EB3",x"B501",x"2F23",x"A00A",x"A009",x"3FFF",x"A008",x"2F23",x"A00A",x"4286", -- 1030-103F
  x"B412",x"B603",x"A007",x"4B7C",x"B434",x"B434",x"B502",x"A00A",x"502C",x"B502",x"A009",x"B434",x"428D",x"B501",x"9005",x"B434", -- 1040-104F
  x"4286",x"B434",x"4286",x"8FF2",x"B200",x"B300",x"8001",x"4D01",x"A003",x"FFCF",x"35A9",x"0004",x"4781",x"B501",x"4EC3",x"9006", -- 1050-105F
  x"4EB3",x"B412",x"B300",x"3FFF",x"A008",x"8002",x"B300",x"0001",x"A003",x"FFF0",x"35AE",x"0005",x"4069",x"2F2B",x"FFFB",x"35B4", -- 1060-106F
  x"0005",x"4069",x"2F2C",x"FFFB",x"35BA",x"0005",x"4069",x"2F2D",x"FFFB",x"35C0",x"0007",x"4781",x"2F2C",x"A00A",x"900F",x"436D", -- 1070-107F
  x"436D",x"35C8",x"0008",x"41F5",x"2F23",x"4366",x"42E2",x"B60C",x"4FA7",x"B603",x"4FA7",x"42CF",x"B501",x"4F88",x"FFFF",x"2D04", -- 1080-108F
  x"A009",x"A003",x"FFE6",x"35D1",x"0007",x"4781",x"0000",x"2D04",x"A009",x"2F2C",x"A00A",x"900B",x"436D",x"436D",x"35D9",x"0008", -- 1090-109F
  x"41F5",x"2F23",x"4366",x"B502",x"4F88",x"B501",x"4F88",x"A003",x"FFEA",x"35E2",x"000C",x"4781",x"0008",x"43FB",x"4C86",x"4415", -- 10A0-10AF
  x"A009",x"507C",x"B502",x"505D",x"441D",x"A009",x"B501",x"505D",x"4426",x"A009",x"444A",x"A009",x"4441",x"A009",x"B412",x"4453", -- 10B0-10BF
  x"A009",x"441D",x"A00A",x"442F",x"A009",x"FFFF",x"442F",x"42C4",x"B502",x"442F",x"A00A",x"4EDD",x"4426",x"A00A",x"4438",x"A009", -- 10C0-10CF
  x"FFFF",x"4438",x"42C4",x"4C86",x"B434",x"B434",x"B412",x"B502",x"4438",x"A00A",x"4EDD",x"B502",x"4D40",x"4441",x"A00A",x"442F", -- 10D0-10DF
  x"A00A",x"4EDD",x"444A",x"A00A",x"4438",x"A00A",x"4EDD",x"4D40",x"4D34",x"4453",x"A00A",x"4D4C",x"B43C",x"B412",x"4C8D",x"B412", -- 10E0-10EF
  x"4D01",x"B412",x"4438",x"A00A",x"B434",x"4F00",x"4438",x"A00A",x"A00D",x"9FD6",x"B434",x"442F",x"A00A",x"B434",x"4F00",x"B412", -- 10F0-10FF
  x"442F",x"A00A",x"A00D",x"9FC1",x"4D01",x"4415",x"A00A",x"4C8D",x"B412",x"4FD9",x"B412",x"4D01",x"FFFF",x"2F2B",x"42C4",x"5096", -- 1100-110F
  x"4409",x"A003",x"FF96",x"35EF",x"000B",x"4781",x"0008",x"43FB",x"4C86",x"4415",x"A009",x"441D",x"A009",x"0001",x"0000",x"4426", -- 1110-111F
  x"A009",x"4453",x"A009",x"0000",x"4441",x"A009",x"0000",x"444A",x"A009",x"B501",x"4426",x"A00A",x"4EDD",x"4426",x"A00A",x"4EDD", -- 1120-112F
  x"441D",x"A00A",x"442F",x"A009",x"FFFF",x"442F",x"42C4",x"B502",x"442F",x"A00A",x"4EDD",x"4426",x"A00A",x"4EDD",x"4441",x"A00A", -- 1130-113F
  x"442F",x"A00A",x"B434",x"4F00",x"4441",x"A009",x"B502",x"4426",x"A00A",x"4EDD",x"442F",x"A00A",x"4EDD",x"444A",x"A00A",x"442F", -- 1140-114F
  x"A00A",x"B434",x"4F00",x"444A",x"A009",x"442F",x"A00A",x"A00D",x"9FDB",x"4441",x"A00A",x"4426",x"A00A",x"4EDD",x"4453",x"A00A", -- 1150-115F
  x"4D28",x"4441",x"A00A",x"4426",x"A00A",x"B434",x"4F00",x"4441",x"A009",x"444A",x"A00A",x"4426",x"A00A",x"4EDD",x"4453",x"A00A", -- 1160-116F
  x"4D34",x"444A",x"A00A",x"4426",x"A00A",x"B434",x"4F00",x"444A",x"A009",x"4453",x"A00A",x"B412",x"4441",x"A00A",x"444A",x"A00A", -- 1170-117F
  x"50AC",x"0001",x"4426",x"42C4",x"4426",x"A00A",x"441D",x"A00A",x"429B",x"9F97",x"4415",x"A00A",x"4C8D",x"B412",x"4FD9",x"B412", -- 1180-118F
  x"4D01",x"4409",x"A003",x"FF7F",x"35FB",x"0011",x"4781",x"0003",x"43FB",x"4415",x"A009",x"0000",x"4415",x"A00A",x"441D",x"A009", -- 1190-119F
  x"441D",x"A00A",x"B501",x"901F",x"428D",x"441D",x"A009",x"441D",x"A00A",x"4EF9",x"4415",x"A00A",x"4426",x"A009",x"4426",x"A00A", -- 11A0-11AF
  x"B501",x"900E",x"428D",x"4426",x"A009",x"4426",x"A00A",x"441D",x"A00A",x"4286",x"4426",x"A00A",x"4286",x"4E42",x"4F00",x"8FEE", -- 11B0-11BF
  x"B300",x"4F00",x"8FDD",x"B300",x"4409",x"A003",x"FFCD",x"360D",x"0005",x"4781",x"2F11",x"A00A",x"B501",x"4286",x"A00A",x"B502", -- 11C0-11CF
  x"0002",x"A007",x"A00A",x"433C",x"0020",x"431D",x"B501",x"A00A",x"9004",x"B501",x"A00A",x"A007",x"8FEF",x"B300",x"A003",x"FFE7", -- 11D0-11DF
  x"3613",x"0005",x"4781",x"2F11",x"A00A",x"B501",x"0004",x"A007",x"435E",x"B501",x"4286",x"A00A",x"B502",x"0002",x"A007",x"A00A", -- 11E0-11EF
  x"433C",x"0020",x"431D",x"B501",x"A00A",x"9004",x"B501",x"A00A",x"A007",x"8FEB",x"B300",x"A003",x"FFE3",x"3619",x"0006",x"4781", -- 11F0-11FF
  x"0020",x"45E4",x"465E",x"900E",x"2F0F",x"A009",x"41FB",x"B501",x"A00A",x"A007",x"2F11",x"A009",x"41FB",x"4286",x"A00A",x"2F13", -- 1200-120F
  x"A009",x"8004",x"B300",x"3620",x"000F",x"41F5",x"A003",x"FFE5",x"3630",x"000A",x"4781",x"436D",x"B501",x"0000",x"429B",x"9003", -- 1210-121F
  x"363B",x"0013",x"41F5",x"B501",x"0003",x"429B",x"9003",x"364F",x"0014",x"41F5",x"B501",x"0006",x"429B",x"9003",x"3664",x"0014", -- 1220-122F
  x"41F5",x"B501",x"0009",x"429B",x"9003",x"3679",x"0030",x"41F5",x"B501",x"0012",x"429B",x"9003",x"36AA",x"0012",x"41F5",x"B501", -- 1230-123F
  x"0369",x"429B",x"9003",x"36BD",x"0013",x"41F5",x"B501",x"1234",x"429B",x"9003",x"36D1",x"0034",x"41F5",x"A003",x"FFC9",x"3706", -- 1240-124F
  x"0005",x"4781",x"47A1",x"41FB",x"0003",x"4294",x"B501",x"435E",x"A00A",x"4286",x"B501",x"435E",x"A00A",x"B501",x"435E",x"0040", -- 1250-125F
  x"4294",x"41FB",x"B412",x"0007",x"A008",x"2F18",x"A007",x"A009",x"A003",x"FFE5",x"370C",x"0002",x"4781",x"0007",x"431D",x"370F", -- 1260-126F
  x"0008",x"41F5",x"A003",x"FFF6",x"3718",x"0002",x"4781",x"0007",x"431D",x"371B",x"0004",x"41F5",x"4713",x"A003",x"FFF5",x"3720", -- 1270-127F
  x"0002",x"4781",x"3723",x"0029",x"41F5",x"436D",x"3A00",x"0100",x"44D2",x"46C6",x"374D",x"0002",x"41F5",x"A003",x"FFF0",x"3750", -- 1280-128F
  x"0005",x"4781",x"2F09",x"A00A",x"0100",x"44D2",x"A003",x"FFF7",x"3756",x"0007",x"4773",x"003C",x"431D",x"375E",x"0004",x"41F5", -- 1290-129F
  x"436D",x"5292",x"3763",x"0007",x"41EF",x"462A",x"9FF9",x"003C",x"431D",x"376B",x"0003",x"41F5",x"A003",x"FFEA",x"376F",x"0003", -- 12A0-12AF
  x"4781",x"0010",x"2F08",x"A009",x"A003",x"FFF8",x"3773",x"0007",x"4781",x"000A",x"2F08",x"A009",x"A003",x"FFF8",x"377B",x"0001", -- 12B0-12BF
  x"4781",x"A00A",x"4F88",x"A003",x"FFF9",x"377D",x"0002",x"4781",x"B501",x"4286",x"A00A",x"B412",x"A00A",x"A003",x"FFF6",x"3780", -- 12C0-12CF
  x"0002",x"4781",x"B412",x"B502",x"A009",x"4286",x"A009",x"A003",x"FFF6",x"3783",x"0002",x"4781",x"52C8",x"4FA7",x"A003",x"FFF9", -- 12D0-12DF
  x"3786",x"0005",x"4069",x"2F2E",x"FFFB",x"378C",x"0006",x"4781",x"A000",x"2F2E",x"42C4",x"2F2E",x"A00A",x"4074",x"A003",x"FFF5", -- 12E0-12EF
  x"3793",x"0006",x"4069",x"2EE0",x"FFFB",x"379A",x"000D",x"4069",x"2F2F",x"FFFB",x"37A8",x"0006",x"4781",x"2EE0",x"2F2F",x"A00A", -- 12F0-12FF
  x"B502",x"42A9",x"900C",x"B501",x"A00A",x"436D",x"B501",x"435E",x"0003",x"4294",x"52C8",x"B412",x"433C",x"4286",x"8FEF",x"B300", -- 1300-130F
  x"A003",x"FFE8",x"37AF",x"0007",x"4069",x"2F30",x"FFFB",x"37B7",x"0008",x"4069",x"2F31",x"FFFB",x"37C0",x"0007",x"4069",x"2F32", -- 1310-131F
  x"FFFB",x"37C8",x"0004",x"4781",x"2F10",x"A00A",x"2F31",x"A009",x"0000",x"2F10",x"A009",x"2EE0",x"B501",x"2F2F",x"A00A",x"42A2", -- 1320-132F
  x"9007",x"B501",x"42E2",x"A00A",x"430B",x"42CF",x"4286",x"8FF4",x"B300",x"2F31",x"A00A",x"2F10",x"A009",x"A003",x"FFE2",x"37CD", -- 1330-133F
  x"0008",x"4781",x"0020",x"45E4",x"465E",x"469E",x"B300",x"4286",x"0000",x"2F30",x"A009",x"2EE0",x"2F2F",x"A00A",x"B502",x"42A9", -- 1340-134F
  x"9014",x"B603",x"A00A",x"429B",x"9006",x"0001",x"2F30",x"A009",x"FFFF",x"2F2F",x"42C4",x"2F30",x"A00A",x"9005",x"B501",x"4286", -- 1350-135F
  x"A00A",x"B502",x"A009",x"4286",x"8FE7",x"B300",x"2F30",x"A009",x"A003",x"FFD5",x"37D6",x"0009",x"4781",x"5342",x"2F30",x"A00A", -- 1360-136F
  x"2F2F",x"A00A",x"A009",x"0001",x"2F2F",x"42C4",x"A003",x"FFF2",x"37E0",x"0011",x"4069",x"2804",x"FFFB",x"37F2",x"0012",x"4069", -- 1370-137F
  x"2804",x"FFFB",x"3805",x"0010",x"4069",x"2805",x"FFFB",x"3816",x"0011",x"4069",x"2805",x"FFFB",x"3828",x"0010",x"4069",x"2806", -- 1380-138F
  x"FFFB",x"3839",x"0011",x"4069",x"2806",x"FFFB",x"384B",x"000F",x"4069",x"2807",x"FFFB",x"385B",x"0010",x"4069",x"2807",x"FFFB", -- 1390-139F
  x"386C",x"000C",x"4781",x"0007",x"0800",x"4047",x"A003",x"FFF8",x"3879",x"000B",x"4781",x"0007",x"0C00",x"4047",x"A003",x"FFF8", -- 13A0-13AF
  x"3885",x"000B",x"4781",x"0007",x"0800",x"4047",x"A003",x"FFF8",x"3891",x"000A",x"4781",x"0007",x"0C00",x"4047",x"A003",x"FFF8", -- 13B0-13BF
  x"389C",x"0005",x"4069",x"2F33",x"FFFB",x"38A2",x"0005",x"4069",x"2F34",x"FFFB",x"38A8",x"0005",x"4069",x"2F35",x"FFFB",x"38AE", -- 13C0-13CF
  x"0005",x"4069",x"2F36",x"FFFB",x"38B4",x"0002",x"4069",x"2F37",x"FFFB",x"38B7",x"0002",x"4069",x"2F38",x"FFFB",x"38BA",x"000A", -- 13D0-13DF
  x"4069",x"2F39",x"FFFB",x"38C5",x"0009",x"4069",x"2F3A",x"FFFB",x"38CF",x"000B",x"4069",x"2F3B",x"FFFB",x"38DB",x"000A",x"4069", -- 13E0-13EF
  x"2F3C",x"FFFB",x"38E6",x"0009",x"4781",x"0001",x"43FB",x"4415",x"A009",x"2F2D",x"A00A",x"9011",x"436D",x"003A",x"431D",x"4415", -- 13F0-13FF
  x"A00A",x"431D",x"0020",x"431D",x"4FA7",x"4415",x"A00A",x"431D",x"003A",x"431D",x"0020",x"431D",x"8001",x"B200",x"4409",x"A003", -- 1400-140F
  x"FFE1",x"38F0",x"000C",x"4781",x"2805",x"A00A",x"2F3B",x"A00A",x"4294",x"9007",x"2F2D",x"A00A",x"9004",x"436D",x"38FD",x"0007", -- 1410-141F
  x"41F5",x"2805",x"A00A",x"2F3B",x"A00A",x"4294",x"9001",x"8FF9",x"53A3",x"A009",x"B501",x"9008",x"B412",x"B502",x"53A3",x"0005", -- 1420-142F
  x"A007",x"B412",x"4851",x"8005",x"B412",x"53A3",x"0005",x"A007",x"A009",x"B501",x"53A3",x"0004",x"A007",x"A009",x"4C86",x"B434", -- 1430-143F
  x"B434",x"53A3",x"0006",x"A007",x"A007",x"2F23",x"A009",x"2F25",x"A00A",x"B412",x"2F27",x"A00A",x"9004",x"0007",x"0C00",x"4047", -- 1440-144F
  x"8001",x"2400",x"2F25",x"A009",x"502C",x"B412",x"2F25",x"A009",x"B412",x"4C8D",x"53A3",x"0003",x"A007",x"A009",x"B603",x"0072", -- 1450-145F
  x"53F5",x"53A3",x"0002",x"A007",x"A009",x"53A3",x"0001",x"A007",x"A009",x"2805",x"A00A",x"A00B",x"0001",x"A008",x"2F3B",x"A009", -- 1460-146F
  x"2805",x"A00A",x"A00B",x"2804",x"A009",x"A003",x"FF9A",x"3905",x"000C",x"4781",x"2807",x"A00A",x"2F3C",x"A00A",x"4294",x"9007", -- 1470-147F
  x"2F2D",x"A00A",x"9004",x"436D",x"3912",x"0007",x"41F5",x"2807",x"A00A",x"2F3C",x"A00A",x"4294",x"9001",x"8FF9",x"53AB",x"A009", -- 1480-148F
  x"B501",x"9008",x"B412",x"B502",x"53AB",x"0005",x"A007",x"B412",x"4851",x"8005",x"B412",x"53AB",x"0005",x"A007",x"A009",x"B501", -- 1490-149F
  x"53AB",x"0004",x"A007",x"A009",x"4C86",x"B434",x"B434",x"53AB",x"0006",x"A007",x"A007",x"2F23",x"A009",x"2F25",x"A00A",x"B412", -- 14A0-14AF
  x"2F27",x"A00A",x"9004",x"0008",x"0000",x"4047",x"8001",x"2800",x"2F25",x"A009",x"502C",x"B412",x"2F25",x"A009",x"B412",x"4C8D", -- 14B0-14BF
  x"53AB",x"0003",x"A007",x"A009",x"B603",x"0075",x"53F5",x"53AB",x"0002",x"A007",x"A009",x"53AB",x"0001",x"A007",x"A009",x"2807", -- 14C0-14CF
  x"A00A",x"A00B",x"0001",x"A008",x"2F3C",x"A009",x"2807",x"A00A",x"A00B",x"2806",x"A009",x"A003",x"FF9A",x"391A",x"000A",x"4781", -- 14D0-14DF
  x"0006",x"43FB",x"4441",x"A009",x"4438",x"A009",x"442F",x"A009",x"4426",x"A009",x"441D",x"A009",x"4415",x"A009",x"4415",x"A00A", -- 14E0-14EF
  x"441D",x"A00A",x"4426",x"A00A",x"442F",x"A00A",x"4438",x"A00A",x"4441",x"A00A",x"4415",x"A00A",x"441D",x"A00A",x"B502",x"902D", -- 14F0-14FF
  x"B200",x"547A",x"4441",x"A00A",x"0003",x"429B",x"441D",x"A00A",x"A00D",x"A00B",x"A008",x"900B",x"0000",x"441D",x"A00A",x"4426", -- 1500-150F
  x"A00A",x"442F",x"A00A",x"4438",x"A00A",x"0002",x"5414",x"4441",x"A00A",x"0003",x"429B",x"9010",x"4426",x"A00A",x"442F",x"A00A", -- 1510-151F
  x"4438",x"A00A",x"B501",x"9002",x"46C6",x"8006",x"B300",x"B501",x"9002",x"430B",x"8001",x"B300",x"802F",x"B501",x"901D",x"B200", -- 1520-152F
  x"5414",x"4441",x"A00A",x"0002",x"429B",x"4441",x"A00A",x"0003",x"429B",x"A00E",x"9010",x"4426",x"A00A",x"442F",x"A00A",x"4438", -- 1530-153F
  x"A00A",x"B501",x"9002",x"46C6",x"8006",x"B300",x"B501",x"9002",x"430B",x"8001",x"B300",x"8010",x"B200",x"B200",x"B43C",x"B200", -- 1540-154F
  x"4438",x"A00A",x"B501",x"9002",x"46C6",x"8006",x"B300",x"B501",x"9002",x"430B",x"8001",x"B300",x"4409",x"A003",x"FF7E",x"3925", -- 1550-155F
  x"0006",x"4781",x"2F2B",x"A00A",x"9002",x"5324",x"8FFB",x"A003",x"FFF6",x"392C",x"0007",x"4781",x"4CB4",x"2F2B",x"A00A",x"A00D", -- 1560-156F
  x"9003",x"FFFF",x"2F2B",x"A009",x"2F2D",x"A00A",x"9009",x"436D",x"3934",x"0003",x"41F5",x"B603",x"4FA7",x"3938",x"0003",x"41F5", -- 1570-157F
  x"B502",x"2F35",x"A00A",x"42A2",x"B502",x"2F36",x"A00A",x"42A2",x"A008",x"900C",x"FFFF",x"2F33",x"A009",x"FFFF",x"2F34",x"A009", -- 1580-158F
  x"FFFF",x"2F35",x"A009",x"FFFF",x"2F36",x"A009",x"B502",x"2F33",x"A00A",x"429B",x"A00B",x"2F35",x"A00A",x"FFFF",x"429B",x"A008", -- 1590-159F
  x"9027",x"2F33",x"A00A",x"FFFF",x"429B",x"9004",x"B502",x"2F33",x"A009",x"800A",x"B502",x"2F35",x"A009",x"2F35",x"A00A",x"2F33", -- 15A0-15AF
  x"A00A",x"4294",x"2F37",x"A009",x"2F2D",x"A00A",x"9009",x"436D",x"2F33",x"4366",x"2F34",x"4366",x"2F35",x"4366",x"2F36",x"4366", -- 15B0-15BF
  x"B502",x"4286",x"B502",x"0000",x"0000",x"0000",x"0000",x"547A",x"B501",x"2F34",x"A00A",x"429B",x"A00B",x"2F36",x"A00A",x"FFFF", -- 15C0-15CF
  x"429B",x"A008",x"9027",x"2F34",x"A00A",x"FFFF",x"429B",x"9004",x"B501",x"2F34",x"A009",x"800A",x"B501",x"2F36",x"A009",x"2F36", -- 15D0-15DF
  x"A00A",x"2F34",x"A00A",x"4294",x"2F38",x"A009",x"2F2D",x"A00A",x"9009",x"436D",x"2F33",x"4366",x"2F34",x"4366",x"2F35",x"4366", -- 15E0-15EF
  x"2F36",x"4366",x"B502",x"B502",x"4286",x"0000",x"0000",x"0000",x"0000",x"5414",x"B200",x"2F35",x"A00A",x"FFFF",x"429B",x"2F36", -- 15F0-15FF
  x"A00A",x"FFFF",x"429B",x"A00E",x"9002",x"5562",x"8003",x"0000",x"2F2B",x"A009",x"A003",x"FF5D",x"393C",x"0008",x"4781",x"0001", -- 1600-160F
  x"43FB",x"4415",x"A009",x"4415",x"A00A",x"0003",x"A007",x"A00A",x"4415",x"A00A",x"0005",x"A007",x"4415",x"A00A",x"0004",x"A007", -- 1610-161F
  x"A00A",x"A00D",x"9001",x"A00A",x"4415",x"A00A",x"0004",x"A007",x"A00A",x"4409",x"A003",x"FFE0",x"3945",x"0008",x"4781",x"0001", -- 1620-162F
  x"43FB",x"4415",x"A009",x"2F2D",x"A00A",x"901C",x"003A",x"431D",x"4415",x"A00A",x"431D",x"0020",x"431D",x"B434",x"B501",x"4F88", -- 1630-163F
  x"B434",x"B434",x"B501",x"9005",x"B603",x"433C",x"0020",x"431D",x"8002",x"B502",x"435E",x"4415",x"A00A",x"431D",x"003A",x"431D", -- 1640-164F
  x"0020",x"431D",x"4409",x"A003",x"FFD7",x"394E",x"0008",x"4781",x"B501",x"9002",x"46C6",x"8006",x"B300",x"B501",x"9002",x"430B", -- 1650-165F
  x"8001",x"B300",x"A003",x"FFF1",x"3957",x"0008",x"4781",x"2F39",x"A00A",x"2804",x"A00A",x"429B",x"A00B",x"9063",x"53B3",x"A00A", -- 1660-166F
  x"A00D",x"9010",x"53B3",x"4286",x"B501",x"A00A",x"B412",x"4286",x"A00A",x"2804",x"A00A",x"2F39",x"A009",x"2804",x"A00A",x"2805", -- 1670-167F
  x"A009",x"556C",x"53B3",x"A00A",x"0001",x"429B",x"53B3",x"A00A",x"0002",x"429B",x"A00E",x"9045",x"53B3",x"0002",x"A007",x"A00A", -- 1680-168F
  x"428D",x"9032",x"53B3",x"4286",x"A00A",x"53B3",x"0002",x"A007",x"A00A",x"428D",x"B603",x"006C",x"53F5",x"53B3",x"560F",x"53B3", -- 1690-169F
  x"A00A",x"2F36",x"A00A",x"0001",x"429B",x"900A",x"2804",x"A00A",x"2F39",x"A009",x"2804",x"A00A",x"2805",x"A009",x"5414",x"8013", -- 16A0-16AF
  x"5414",x"53B3",x"A00A",x"0002",x"429B",x"9005",x"53B3",x"560F",x"006D",x"562F",x"5658",x"2804",x"A00A",x"2F39",x"A009",x"2804", -- 16B0-16BF
  x"A00A",x"2805",x"A009",x"800D",x"53B3",x"560F",x"006E",x"562F",x"5658",x"2804",x"A00A",x"2F39",x"A009",x"2804",x"A00A",x"2805", -- 16C0-16CF
  x"A009",x"A003",x"FF91",x"3960",x"0008",x"4781",x"2F3A",x"A00A",x"2806",x"A00A",x"429B",x"A00B",x"90A2",x"53BB",x"A00A",x"A00D", -- 16D0-16DF
  x"9010",x"53BB",x"4286",x"B501",x"A00A",x"B412",x"4286",x"A00A",x"2806",x"A00A",x"2F3A",x"A009",x"2806",x"A00A",x"2807",x"A009", -- 16E0-16EF
  x"556C",x"53BB",x"A00A",x"0001",x"429B",x"53BB",x"A00A",x"0003",x"429B",x"A00E",x"9084",x"53BB",x"4286",x"A00A",x"428D",x"9044", -- 16F0-16FF
  x"53BB",x"4286",x"A00A",x"428D",x"53BB",x"0002",x"A007",x"A00A",x"B603",x"006F",x"53F5",x"53BB",x"560F",x"53BB",x"A00A",x"2F35", -- 1700-170F
  x"A00A",x"0001",x"429B",x"900A",x"2806",x"A00A",x"2F3A",x"A009",x"2806",x"A00A",x"2807",x"A009",x"547A",x"8025",x"547A",x"53BB", -- 1710-171F
  x"A00A",x"0003",x"429B",x"9017",x"53BB",x"0002",x"A007",x"A00A",x"900D",x"0000",x"53BB",x"0002",x"A007",x"A00A",x"53BB",x"560F", -- 1720-172F
  x"B434",x"502C",x"B434",x"B434",x"0002",x"5414",x"53BB",x"560F",x"004D",x"562F",x"5658",x"2806",x"A00A",x"2F3A",x"A009",x"2806", -- 1730-173F
  x"A00A",x"2807",x"A009",x"803B",x"53BB",x"0002",x"A007",x"A00A",x"9029",x"53BB",x"4286",x"A00A",x"428D",x"53BB",x"0002",x"A007", -- 1740-174F
  x"A00A",x"B603",x"004F",x"53F5",x"53BB",x"560F",x"B434",x"502C",x"B434",x"B434",x"53BB",x"A00A",x"0003",x"429B",x"9008",x"0002", -- 1750-175F
  x"5414",x"53BB",x"560F",x"004B",x"562F",x"5658",x"8002",x"0001",x"5414",x"2806",x"A00A",x"2F3A",x"A009",x"2806",x"A00A",x"2807", -- 1760-176F
  x"A009",x"800D",x"53BB",x"560F",x"004E",x"562F",x"5658",x"2806",x"A00A",x"2F3A",x"A009",x"2806",x"A00A",x"2807",x"A009",x"A003", -- 1770-177F
  x"FF52",x"3969",x"0001",x"4069",x"2F3D",x"FFFB",x"396B",x"0002",x"4069",x"2F3E",x"FFFB",x"396E",x"0002",x"4069",x"2F3F",x"FFFB", -- 1780-178F
  x"3971",x"0004",x"4069",x"2F40",x"FFFB",x"3976",x"0004",x"4069",x"2F41",x"FFFB",x"397B",x"0006",x"4069",x"2F42",x"FFFB",x"3982", -- 1790-179F
  x"0002",x"4781",x"49E2",x"B412",x"B300",x"A003",x"FFF8",x"3985",x"0005",x"4781",x"2F40",x"A009",x"A003",x"FFF9",x"398B",x"0005", -- 17A0-17AF
  x"4781",x"2F41",x"A009",x"A003",x"FFF9",x"3991",x"0004",x"4781",x"0003",x"43FB",x"B502",x"505D",x"441D",x"A009",x"4426",x"A009", -- 17B0-17BF
  x"4415",x"A009",x"0000",x"441D",x"A00A",x"428D",x"B501",x"441D",x"A009",x"4415",x"A00A",x"B502",x"4EDD",x"4426",x"A00A",x"4EDD", -- 17C0-17CF
  x"4F00",x"441D",x"A00A",x"B501",x"A00D",x"9FEF",x"B300",x"4409",x"A003",x"FFDB",x"3996",x"0005",x"4069",x"2F43",x"FFFB",x"399C", -- 17D0-17DF
  x"0006",x"4069",x"2F44",x"FFFB",x"39A3",x"0004",x"4069",x"2F45",x"FFFB",x"39A8",x"0005",x"4069",x"2F46",x"FFFB",x"39AE",x"0004", -- 17E0-17EF
  x"4781",x"2F44",x"A00A",x"B501",x"0000",x"4EDD",x"B412",x"0001",x"4EDD",x"2F46",x"A00A",x"50AC",x"B412",x"502C",x"B412",x"4D01", -- 17F0-17FF
  x"4CB4",x"B412",x"502C",x"B412",x"4D01",x"A003",x"FFE7",x"39B3",x"0008",x"4781",x"502C",x"2F44",x"A009",x"FFFF",x"2F43",x"A009", -- 1800-180F
  x"2F43",x"A00A",x"2F45",x"A00A",x"A008",x"900D",x"57F1",x"0000",x"2F43",x"A009",x"0000",x"2F45",x"A009",x"0000",x"2F44",x"A009", -- 1810-181F
  x"0000",x"2F46",x"A009",x"A003",x"FFE2",x"39BC",x"0007",x"4781",x"502C",x"2F46",x"A009",x"FFFF",x"2F45",x"A009",x"2F43",x"A00A", -- 1820-182F
  x"2F45",x"A00A",x"A008",x"900D",x"57F1",x"0000",x"2F43",x"A009",x"0000",x"2F45",x"A009",x"0000",x"2F44",x"A009",x"0000",x"2F46", -- 1830-183F
  x"A009",x"A003",x"B501",x"2F0E",x"A009",x"4CB4",x"2F33",x"A00A",x"2F34",x"A00A",x"A00E",x"901F",x"2F33",x"A00A",x"9007",x"2F37", -- 1840-184F
  x"A00A",x"428D",x"2F33",x"A00A",x"4D34",x"8001",x"0000",x"2F34",x"A00A",x"9007",x"2F38",x"A00A",x"428D",x"2F34",x"A00A",x"4D34", -- 1850-185F
  x"8001",x"0000",x"2F0E",x"A00A",x"39C4",x"0012",x"41EF",x"0003",x"54E0",x"8FFF",x"801A",x"0000",x"2F10",x"A009",x"436D",x"2F0A", -- 1860-186F
  x"A00A",x"2F0C",x"A00A",x"2F0A",x"A00A",x"4294",x"428D",x"433C",x"39D7",x"0003",x"41F5",x"39DB",x"000A",x"41EF",x"46C6",x"436D", -- 1870-187F
  x"39E6",x"0016",x"41F5",x"435E",x"8FFF",x"A003",x"FF9E",x"39FD",x"0004",x"4781",x"2F2D",x"A00A",x"9008",x"3A02",x"0005",x"41F5", -- 1880-188F
  x"B603",x"4FA7",x"2F44",x"A00A",x"4F88",x"B502",x"2F40",x"A00A",x"4EDD",x"502C",x"2F2D",x"A00A",x"9002",x"B501",x"4F88",x"2F37", -- 1890-189F
  x"A00A",x"428D",x"0000",x"B434",x"2F33",x"A00A",x"2F34",x"A00A",x"429B",x"9008",x"502C",x"2F41",x"A00A",x"4EF9",x"2F42",x"A00A", -- 18A0-18AF
  x"4D34",x"4F00",x"2F2D",x"A00A",x"9002",x"B501",x"4F88",x"1828",x"0000",x"0003",x"54E0",x"A003",x"FFCA",x"3A08",x"0005",x"4781", -- 18B0-18BF
  x"0005",x"43FB",x"2F2D",x"A00A",x"9005",x"3A0E",x"0006",x"41F5",x"B501",x"4F88",x"2F41",x"A00A",x"B60C",x"B300",x"B412",x"57B8", -- 18C0-18CF
  x"2F2D",x"A00A",x"9002",x"B501",x"4F88",x"0000",x"2F38",x"A00A",x"428D",x"B434",x"2F33",x"A00A",x"2F34",x"A00A",x"429B",x"9008", -- 18D0-18DF
  x"502C",x"2F40",x"A00A",x"4EF9",x"2F42",x"A00A",x"4D28",x"4F00",x"180A",x"2F2D",x"A00A",x"9002",x"B502",x"4F88",x"4438",x"A009", -- 18E0-18EF
  x"442F",x"A009",x"4426",x"A009",x"441D",x"A009",x"4415",x"A009",x"441D",x"A00A",x"4426",x"A00A",x"4FB4",x"4415",x"A00A",x"442F", -- 18F0-18FF
  x"A00A",x"4FBF",x"4438",x"A00A",x"0000",x"0002",x"54E0",x"2F33",x"A00A",x"2F34",x"A00A",x"429B",x"900A",x"0000",x"2F38",x"A00A", -- 1900-190F
  x"428D",x"0000",x"3A15",x"000A",x"41EF",x"0002",x"54E0",x"4409",x"A003",x"FFA3",x"3A20",x"0004",x"4781",x"2F2D",x"A00A",x"9003", -- 1910-191F
  x"3A25",x"0005",x"41F5",x"B501",x"2F2B",x"A009",x"2F3E",x"A009",x"B501",x"2F42",x"A009",x"2F3D",x"A00A",x"2F3E",x"A00A",x"4294", -- 1920-192F
  x"2F3F",x"A009",x"0000",x"2F38",x"A00A",x"428D",x"2F3F",x"A00A",x"2F37",x"A00A",x"57A2",x"17AA",x"0000",x"0002",x"54E0",x"2F37", -- 1930-193F
  x"A00A",x"428D",x"0000",x"2F3F",x"A00A",x"2F38",x"A00A",x"57A2",x"17B1",x"0000",x"0003",x"54E0",x"B502",x"2F40",x"A00A",x"4EDD", -- 1940-194F
  x"2F41",x"A00A",x"4EDD",x"2F2D",x"A00A",x"9002",x"B501",x"4F88",x"2F37",x"A00A",x"428D",x"0000",x"B434",x"18C0",x"0000",x"0003", -- 1950-195F
  x"54E0",x"2F3E",x"A00A",x"428D",x"9009",x"0001",x"0001",x"2F3D",x"A00A",x"3A2B",x"0004",x"41EF",x"0001",x"54E0",x"2F3E",x"A00A", -- 1960-196F
  x"428D",x"900A",x"0001",x"0001",x"2F3E",x"A00A",x"428D",x"3A30",x"0005",x"41EF",x"0001",x"54E0",x"A003",x"FF9C",x"3A36",x"0009", -- 1970-197F
  x"4781",x"0007",x"43FB",x"441D",x"A009",x"4415",x"A009",x"2F37",x"A00A",x"428D",x"2F38",x"A00A",x"428D",x"0000",x"3A40",x"0009", -- 1980-198F
  x"41EF",x"0003",x"54E0",x"0000",x"4426",x"A009",x"0000",x"4438",x"A009",x"4415",x"A00A",x"4438",x"A00A",x"4EDD",x"444A",x"A009", -- 1990-199F
  x"0000",x"442F",x"A009",x"0000",x"4441",x"A009",x"4426",x"A00A",x"442F",x"A00A",x"444A",x"A00A",x"4441",x"A00A",x"4EDD",x"0D01", -- 19A0-19AF
  x"0000",x"0001",x"54E0",x"0001",x"442F",x"42C4",x"442F",x"A00A",x"2F38",x"A00A",x"429B",x"9003",x"0000",x"442F",x"A009",x"0001", -- 19B0-19BF
  x"4441",x"42C4",x"4441",x"A00A",x"2F3D",x"A00A",x"429B",x"9FDE",x"0001",x"4426",x"42C4",x"4426",x"A00A",x"2F37",x"A00A",x"429B", -- 19C0-19CF
  x"900F",x"0000",x"4426",x"A009",x"2F37",x"A00A",x"428D",x"2F38",x"A00A",x"428D",x"0000",x"3A4A",x"0009",x"41EF",x"0003",x"54E0", -- 19D0-19DF
  x"0001",x"4438",x"42C4",x"4438",x"A00A",x"2F3D",x"A00A",x"429B",x"9FB0",x"2F37",x"A00A",x"428D",x"2F38",x"A00A",x"428D",x"0000", -- 19E0-19EF
  x"3A54",x"0009",x"41EF",x"0003",x"54E0",x"2F37",x"A00A",x"428D",x"2F38",x"A00A",x"428D",x"441D",x"A00A",x"0000",x"0000",x"0003", -- 19F0-19FF
  x"54E0",x"4409",x"A003",x"FF7A",x"3A5E",x"0012",x"4781",x"2F3D",x"A00A",x"591D",x"5562",x"A003",x"FFF7",x"3A71",x"0005",x"4781", -- 1A00-1A0F
  x"2F2D",x"A00A",x"9003",x"3A77",x"0006",x"41F5",x"0001",x"2F2B",x"A009",x"0001",x"2F3E",x"A009",x"2F42",x"A009",x"0000",x"2F38", -- 1A10-1A1F
  x"A00A",x"428D",x"0000",x"17AA",x"0000",x"0002",x"54E0",x"2F37",x"A00A",x"428D",x"0000",x"0000",x"17B1",x"0000",x"0003",x"54E0", -- 1A20-1A2F
  x"B502",x"2F40",x"A00A",x"4EDD",x"2F41",x"A00A",x"4EDD",x"B501",x"4F88",x"2F42",x"A00A",x"4D40",x"B502",x"4D28",x"B501",x"4F88", -- 1A30-1A3F
  x"0000",x"2F42",x"A009",x"2F37",x"A00A",x"428D",x"0000",x"B434",x"18C0",x"0000",x"0003",x"54E0",x"5562",x"A003",x"FFBE",x"3A7E", -- 1A40-1A4F
  x"0007",x"4781",x"0000",x"2F2B",x"A009",x"A003",x"FFF8",x"3A86",x"000F",x"4781",x"0001",x"43FB",x"4415",x"A009",x"B502",x"4415", -- 1A50-1A5F
  x"A00A",x"0000",x"4EDD",x"4EDD",x"4415",x"A00A",x"0001",x"4EDD",x"4EDD",x"2F33",x"A00A",x"9006",x"2F37",x"A00A",x"2F33",x"A00A", -- 1A60-1A6F
  x"4D34",x"8001",x"0000",x"2F34",x"A00A",x"9006",x"2F38",x"A00A",x"2F34",x"A00A",x"4D34",x"8001",x"0000",x"B434",x"1A52",x"0000", -- 1A70-1A7F
  x"0001",x"54E0",x"4409",x"A003",x"FFD2",x"3A96",x"0007",x"4781",x"0004",x"43FB",x"441D",x"A009",x"4415",x"A009",x"4415",x"A00A", -- 1A80-1A8F
  x"2F37",x"A00A",x"49E2",x"4426",x"A009",x"441D",x"A00A",x"2F38",x"A00A",x"49E2",x"442F",x"A009",x"0001",x"2F2B",x"A009",x"4FB4", -- 1A90-1A9F
  x"4426",x"A00A",x"442F",x"A00A",x"4FBF",x"1A5A",x"0000",x"0001",x"54E0",x"5562",x"4409",x"A003",x"FFD8",x"3A9E",x"0019",x"4781", -- 1AA0-1AAF
  x"2F37",x"A00A",x"428D",x"2F38",x"A00A",x"428D",x"0000",x"0CB4",x"0000",x"0003",x"54E0",x"A003",x"FFF0",x"3AB8",x"000B",x"4781", -- 1AB0-1ABF
  x"2F37",x"A00A",x"428D",x"2F38",x"A00A",x"428D",x"B434",x"0000",x"0000",x"0003",x"54E0",x"A003",x"FFF0",x"3AC4",x"0004",x"4781", -- 1AC0-1ACF
  x"0003",x"43FB",x"4426",x"A009",x"441D",x"A009",x"4415",x"A009",x"441D",x"A00A",x"4EF9",x"4426",x"A00A",x"4415",x"A00A",x"4D01", -- 1AD0-1ADF
  x"4F00",x"4F00",x"4409",x"A003",x"FFE8",x"3AC9",x"0007",x"4781",x"0007",x"43FB",x"4426",x"A009",x"441D",x"A009",x"4415",x"A009", -- 1AE0-1AEF
  x"441D",x"A00A",x"2F37",x"A00A",x"49E2",x"4441",x"A009",x"442F",x"A009",x"4426",x"A00A",x"2F38",x"A00A",x"49E2",x"444A",x"A009", -- 1AF0-1AFF
  x"4438",x"A009",x"442F",x"A00A",x"4438",x"A00A",x"4415",x"A00A",x"0000",x"0000",x"0001",x"54E0",x"442F",x"A00A",x"4438",x"A00A", -- 1B00-1B0F
  x"4441",x"A00A",x"0000",x"0000",x"0001",x"54E0",x"442F",x"A00A",x"4438",x"A00A",x"444A",x"A00A",x"1AD0",x"0000",x"0001",x"54E0", -- 1B10-1B1F
  x"4409",x"A003",x"FFC2",x"3AD1",x"0022",x"4781",x"0003",x"43FB",x"2F3D",x"A009",x"2F3D",x"A00A",x"441D",x"A009",x"441D",x"A00A", -- 1B20-1B2F
  x"B501",x"9028",x"428D",x"441D",x"A009",x"2F3D",x"A00A",x"4426",x"A009",x"4426",x"A00A",x"B501",x"901B",x"428D",x"4426",x"A009", -- 1B30-1B3F
  x"441D",x"A00A",x"4286",x"4426",x"A00A",x"4286",x"4E42",x"2F2D",x"A00A",x"9008",x"436D",x"441D",x"A00A",x"4426",x"A00A",x"4FA7", -- 1B40-1B4F
  x"B501",x"4F88",x"441D",x"A00A",x"4426",x"A00A",x"5AE8",x"8FE1",x"B300",x"8FD4",x"B300",x"4409",x"A003",x"0000",x"0000",x"0000", -- 1B50-1B5F

  SHA(10*16-1 downto 9*16),
  SHA(9*16-1 downto 8*16),
  SHA(8*16-1 downto 7*16),
  SHA(7*16-1 downto 6*16),
  SHA(6*16-1 downto 5*16),
  SHA(5*16-1 downto 4*16),
  SHA(4*16-1 downto 3*16),
  SHA(3*16-1 downto 2*16),
  SHA(2*16-1 downto 1*16),
  SHA(1*16-1 downto 0*16),
  others=>x"0000");

-- Textspeicher
type ByteRAMTYPE is array(0 to 4*1024-1) of STD_LOGIC_VECTOR (7 downto 0);
signal ByteRAM: ByteRAMTYPE:=(

  x"28",x"20",x"7B",x"20",x"7D",x"20",x"43",x"4F",x"4D",x"50",x"49",x"4C",x"45",x"20",x"4D",x"4C", -- 3000-300F
  x"49",x"54",x"20",x"41",x"42",x"53",x"20",x"4C",x"49",x"54",x"2C",x"20",x"28",x"43",x"4F",x"4E", -- 3010-301F
  x"53",x"54",x"41",x"4E",x"54",x"3A",x"29",x"20",x"43",x"4F",x"4E",x"53",x"54",x"41",x"4E",x"54", -- 3020-302F
  x"20",x"4B",x"45",x"59",x"41",x"44",x"52",x"20",x"53",x"50",x"20",x"52",x"50",x"20",x"50",x"43", -- 3030-303F
  x"20",x"58",x"42",x"49",x"54",x"20",x"53",x"4D",x"55",x"44",x"47",x"45",x"42",x"49",x"54",x"20", -- 3040-304F
  x"52",x"50",x"30",x"20",x"49",x"52",x"41",x"4D",x"41",x"44",x"52",x"20",x"4A",x"52",x"41",x"4D", -- 3050-305F
  x"41",x"44",x"52",x"20",x"58",x"4F",x"46",x"46",x"20",x"43",x"52",x"42",x"5A",x"45",x"49",x"47", -- 3060-306F
  x"20",x"43",x"52",x"44",x"50",x"20",x"42",x"41",x"53",x"45",x"20",x"54",x"49",x"42",x"20",x"49", -- 3070-307F
  x"4E",x"31",x"20",x"49",x"4E",x"32",x"20",x"49",x"4E",x"33",x"20",x"49",x"4E",x"34",x"20",x"45", -- 3080-308F
  x"52",x"52",x"4F",x"52",x"4E",x"52",x"20",x"44",x"50",x"20",x"53",x"54",x"41",x"54",x"20",x"4C", -- 3090-309F
  x"46",x"41",x"20",x"42",x"41",x"4E",x"46",x"20",x"42",x"5A",x"45",x"49",x"47",x"20",x"44",x"50", -- 30A0-30AF
  x"4D",x"45",x"52",x"4B",x"20",x"43",x"53",x"50",x"20",x"44",x"55",x"42",x"49",x"54",x"20",x"4C", -- 30B0-30BF
  x"4F",x"43",x"41",x"4C",x"41",x"44",x"52",x"45",x"53",x"53",x"45",x"20",x"56",x"45",x"52",x"53", -- 30C0-30CF
  x"49",x"4F",x"4E",x"20",x"52",x"45",x"54",x"55",x"52",x"4E",x"20",x"28",x"4D",x"43",x"4F",x"44", -- 30D0-30DF
  x"45",x"3A",x"29",x"20",x"4D",x"43",x"4F",x"44",x"45",x"20",x"4D",x"49",x"4E",x"55",x"53",x"20", -- 30E0-30EF
  x"55",x"2B",x"20",x"55",x"2A",x"20",x"30",x"3D",x"20",x"30",x"4C",x"54",x"20",x"45",x"4D",x"49", -- 30F0-30FF
  x"54",x"43",x"4F",x"44",x"45",x"20",x"4E",x"4F",x"54",x"20",x"41",x"4E",x"44",x"20",x"4F",x"52", -- 3100-310F
  x"20",x"4D",x"2B",x"20",x"21",x"20",x"40",x"20",x"53",x"57",x"41",x"50",x"20",x"4F",x"56",x"45", -- 3110-311F
  x"52",x"20",x"44",x"55",x"50",x"20",x"52",x"4F",x"54",x"20",x"44",x"52",x"4F",x"50",x"20",x"32", -- 3120-312F
  x"53",x"57",x"41",x"50",x"20",x"32",x"4F",x"56",x"45",x"52",x"20",x"32",x"44",x"55",x"50",x"20", -- 3130-313F
  x"32",x"44",x"52",x"4F",x"50",x"20",x"4E",x"4F",x"4F",x"50",x"20",x"42",x"2C",x"20",x"5A",x"2C", -- 3140-314F
  x"20",x"28",x"57",x"4F",x"52",x"44",x"3A",x"29",x"20",x"57",x"4F",x"52",x"44",x"3A",x"20",x"22", -- 3150-315F
  x"20",x"2E",x"22",x"20",x"48",x"45",x"52",x"45",x"20",x"4A",x"52",x"42",x"49",x"54",x"20",x"4A", -- 3160-316F
  x"52",x"30",x"42",x"49",x"54",x"20",x"58",x"53",x"45",x"54",x"42",x"54",x"20",x"41",x"4C",x"4C", -- 3170-317F
  x"4F",x"54",x"20",x"42",x"52",x"41",x"4E",x"43",x"48",x"2C",x"20",x"30",x"42",x"52",x"41",x"4E", -- 3180-318F
  x"43",x"48",x"2C",x"20",x"42",x"45",x"47",x"49",x"4E",x"20",x"41",x"47",x"41",x"49",x"4E",x"20", -- 3190-319F
  x"55",x"4E",x"54",x"49",x"4C",x"20",x"49",x"46",x"20",x"45",x"4E",x"44",x"5F",x"49",x"46",x"20", -- 31A0-31AF
  x"45",x"4C",x"53",x"45",x"20",x"57",x"48",x"49",x"4C",x"45",x"20",x"52",x"45",x"50",x"45",x"41", -- 31B0-31BF
  x"54",x"20",x"43",x"40",x"20",x"43",x"21",x"20",x"31",x"2B",x"20",x"31",x"2D",x"20",x"4D",x"2D", -- 31C0-31CF
  x"20",x"3D",x"20",x"4C",x"54",x"20",x"3E",x"20",x"4D",x"2A",x"20",x"42",x"59",x"45",x"20",x"42", -- 31D0-31DF
  x"59",x"45",x"20",x"20",x"2B",x"21",x"20",x"52",x"3E",x"20",x"3E",x"52",x"20",x"52",x"20",x"2C", -- 31E0-31EF
  x"20",x"45",x"58",x"45",x"43",x"55",x"54",x"45",x"20",x"4B",x"45",x"59",x"20",x"45",x"4D",x"49", -- 31F0-31FF
  x"54",x"20",x"53",x"48",x"4C",x"31",x"36",x"20",x"44",x"49",x"47",x"20",x"54",x"59",x"50",x"45", -- 3200-320F
  x"20",x"48",x"47",x"2E",x"20",x"4D",x"2E",x"20",x"4D",x"3F",x"20",x"43",x"52",x"20",x"66",x"6C", -- 3210-321F
  x"3E",x"20",x"2F",x"66",x"6C",x"3E",x"20",x"66",x"72",x"3E",x"20",x"2F",x"66",x"72",x"3E",x"20", -- 3220-322F
  x"46",x"45",x"48",x"4C",x"45",x"52",x"54",x"45",x"58",x"54",x"20",x"44",x"49",x"53",x"41",x"42", -- 3230-323F
  x"4C",x"45",x"20",x"77",x"65",x"69",x"74",x"65",x"72",x"20",x"6E",x"61",x"63",x"68",x"20",x"54", -- 3240-324F
  x"61",x"73",x"74",x"65",x"20",x"45",x"53",x"43",x"41",x"50",x"45",x"20",x"20",x"45",x"52",x"52", -- 3250-325F
  x"4F",x"52",x"20",x"3F",x"3F",x"3F",x"20",x"46",x"45",x"48",x"4C",x"45",x"52",x"54",x"45",x"58", -- 3260-326F
  x"54",x"20",x"45",x"52",x"52",x"4F",x"52",x"20",x"2D",x"20",x"46",x"65",x"68",x"6C",x"65",x"72", -- 3270-327F
  x"20",x"4E",x"75",x"6D",x"6D",x"65",x"72",x"20",x"20",x"43",x"53",x"50",x"21",x"20",x"43",x"53", -- 3280-328F
  x"50",x"3F",x"20",x"4C",x"4F",x"43",x"41",x"4C",x"20",x"45",x"4E",x"44",x"5F",x"4C",x"4F",x"43", -- 3290-329F
  x"41",x"4C",x"20",x"4C",x"30",x"20",x"4C",x"31",x"20",x"4C",x"32",x"20",x"4C",x"33",x"20",x"4C", -- 32A0-32AF
  x"34",x"20",x"4C",x"35",x"20",x"4C",x"36",x"20",x"4C",x"37",x"20",x"27",x"20",x"49",x"4E",x"43", -- 32B0-32BF
  x"52",x"34",x"20",x"4B",x"45",x"59",x"5F",x"49",x"4E",x"54",x"20",x"4B",x"45",x"59",x"43",x"4F", -- 32C0-32CF
  x"44",x"45",x"32",x"20",x"45",x"58",x"50",x"45",x"43",x"54",x"20",x"44",x"49",x"47",x"49",x"54", -- 32D0-32DF
  x"20",x"4E",x"55",x"4D",x"42",x"45",x"52",x"20",x"57",x"4F",x"52",x"44",x"20",x"5A",x"3D",x"20", -- 32E0-32EF
  x"46",x"49",x"4E",x"44",x"20",x"4C",x"43",x"46",x"41",x"20",x"43",x"4F",x"4D",x"50",x"49",x"4C", -- 32F0-32FF
  x"45",x"2C",x"20",x"43",x"52",x"45",x"41",x"54",x"45",x"20",x"49",x"4E",x"54",x"45",x"52",x"50", -- 3300-330F
  x"52",x"45",x"54",x"20",x"51",x"55",x"49",x"54",x"20",x"2F",x"6F",x"6B",x"3E",x"20",x"6F",x"6B", -- 3310-331F
  x"20",x"6F",x"6B",x"3E",x"20",x"2F",x"6F",x"6B",x"3E",x"20",x"6F",x"6B",x"20",x"53",x"54",x"41", -- 3320-332F
  x"52",x"54",x"20",x"46",x"4F",x"52",x"54",x"59",x"2D",x"46",x"4F",x"52",x"54",x"48",x"20",x"53", -- 3330-333F
  x"4D",x"55",x"44",x"47",x"45",x"20",x"28",x"49",x"4D",x"4D",x"45",x"44",x"49",x"41",x"54",x"45", -- 3340-334F
  x"3A",x"29",x"20",x"28",x"43",x"4F",x"4D",x"50",x"49",x"4C",x"45",x"3A",x"29",x"20",x"28",x"3A", -- 3350-335F
  x"29",x"20",x"49",x"4D",x"4D",x"45",x"44",x"49",x"41",x"54",x"45",x"3A",x"20",x"43",x"4F",x"4D", -- 3360-336F
  x"50",x"49",x"4C",x"45",x"3A",x"20",x"3A",x"20",x"3B",x"20",x"4C",x"47",x"2E",x"20",x"4E",x"47", -- 3370-337F
  x"2E",x"20",x"78",x"20",x"2C",x"20",x"44",x"55",x"4D",x"50",x"5A",x"20",x"27",x"20",x"53",x"54", -- 3380-338F
  x"41",x"52",x"54",x"20",x"20",x"44",x"55",x"4D",x"50",x"5A",x"3E",x"20",x"20",x"20",x"20",x"20", -- 3390-339F
  x"2D",x"2D",x"20",x"20",x"2D",x"20",x"2F",x"44",x"55",x"4D",x"50",x"5A",x"3E",x"20",x"52",x"41", -- 33A0-33AF
  x"4D",x"50",x"31",x"20",x"56",x"41",x"52",x"49",x"41",x"42",x"4C",x"45",x"20",x"4D",x"4F",x"56", -- 33B0-33BF
  x"45",x"20",x"46",x"49",x"4C",x"4C",x"20",x"44",x"55",x"4D",x"50",x"20",x"4D",x"41",x"58",x"20", -- 33C0-33CF
  x"4D",x"49",x"4E",x"20",x"4D",x"55",x"4C",x"54",x"5F",x"49",x"20",x"4D",x"55",x"4C",x"54",x"5F", -- 33D0-33DF
  x"49",x"49",x"20",x"53",x"55",x"50",x"45",x"52",x"4D",x"55",x"4C",x"54",x"20",x"41",x"20",x"42", -- 33E0-33EF
  x"20",x"43",x"20",x"53",x"4D",x"55",x"4C",x"20",x"41",x"44",x"44",x"49",x"45",x"52",x"20",x"44", -- 33F0-33FF
  x"49",x"33",x"32",x"20",x"44",x"49",x"56",x"33",x"32",x"20",x"4D",x"2F",x"4D",x"4F",x"44",x"20", -- 3400-340F
  x"53",x"44",x"49",x"56",x"20",x"4F",x"50",x"45",x"52",x"41",x"4E",x"44",x"31",x"20",x"4F",x"50", -- 3410-341F
  x"45",x"52",x"41",x"4E",x"44",x"32",x"20",x"45",x"52",x"47",x"45",x"42",x"4E",x"49",x"53",x"20", -- 3420-342F
  x"5A",x"41",x"48",x"4C",x"45",x"4E",x"53",x"50",x"45",x"49",x"43",x"48",x"45",x"52",x"20",x"53", -- 3430-343F
  x"50",x"45",x"49",x"43",x"48",x"45",x"52",x"45",x"4E",x"44",x"45",x"20",x"53",x"43",x"48",x"49", -- 3440-344F
  x"45",x"42",x"20",x"55",x"42",x"49",x"54",x"20",x"54",x"52",x"49",x"4D",x"20",x"53",x"4C",x"58", -- 3450-345F
  x"2D",x"3E",x"45",x"52",x"47",x"45",x"42",x"4E",x"49",x"53",x"5F",x"4B",x"55",x"52",x"5A",x"20", -- 3460-346F
  x"53",x"4C",x"58",x"2D",x"3E",x"45",x"52",x"47",x"45",x"42",x"4E",x"49",x"53",x"20",x"4F",x"50", -- 3470-347F
  x"45",x"52",x"41",x"4E",x"44",x"2D",x"3E",x"53",x"4C",x"58",x"20",x"45",x"52",x"47",x"45",x"42", -- 3480-348F
  x"4E",x"49",x"53",x"5F",x"4E",x"45",x"55",x"21",x"20",x"49",x"4E",x"49",x"54",x"20",x"53",x"50", -- 3490-349F
  x"45",x"49",x"43",x"48",x"45",x"52",x"48",x"4F",x"4C",x"20",x"32",x"4F",x"50",x"45",x"52",x"41", -- 34A0-34AF
  x"4E",x"44",x"45",x"4E",x"2D",x"3E",x"32",x"53",x"4C",x"58",x"20",x"2B",x"20",x"2D",x"20",x"2A", -- 34B0-34BF
  x"20",x"52",x"45",x"43",x"55",x"52",x"53",x"45",x"20",x"2F",x"4D",x"4F",x"44",x"20",x"48",x"47", -- 34C0-34CF
  x"30",x"2E",x"20",x"2E",x"20",x"2D",x"20",x"42",x"2E",x"20",x"42",x"4C",x"4F",x"43",x"4B",x"41", -- 34D0-34DF
  x"4E",x"46",x"41",x"4E",x"47",x"20",x"42",x"4C",x"4F",x"43",x"4B",x"45",x"4E",x"44",x"45",x"20", -- 34E0-34EF
  x"4E",x"45",x"42",x"45",x"4E",x"52",x"45",x"43",x"48",x"4E",x"55",x"4E",x"47",x"20",x"48",x"41", -- 34F0-34FF
  x"55",x"50",x"54",x"52",x"45",x"43",x"48",x"4E",x"55",x"4E",x"47",x"20",x"52",x"45",x"43",x"48", -- 3500-350F
  x"45",x"4E",x"42",x"4C",x"4F",x"43",x"4B",x"20",x"53",x"50",x"45",x"49",x"43",x"48",x"45",x"52", -- 3510-351F
  x"44",x"41",x"20",x"49",x"4E",x"49",x"54",x"20",x"41",x"2B",x"30",x"20",x"42",x"2B",x"30",x"20", -- 3520-352F
  x"2B",x"20",x"2D",x"20",x"2A",x"20",x"2F",x"20",x"4D",x"4F",x"44",x"20",x"47",x"47",x"54",x"20", -- 3530-353F
  x"42",x"4B",x"20",x"4E",x"4E",x"55",x"4D",x"42",x"45",x"52",x"20",x"4E",x"22",x"20",x"52",x"45", -- 3540-354F
  x"50",x"4C",x"41",x"43",x"45",x"3A",x"20",x"5E",x"20",x"2E",x"20",x"2D",x"20",x"30",x"20",x"20", -- 3550-355F
  x"42",x"2E",x"20",x"5A",x"45",x"52",x"4C",x"45",x"47",x"20",x"4F",x"42",x"4A",x"3F",x"20",x"4C", -- 3560-356F
  x"20",x"47",x"20",x"48",x"20",x"2E",x"20",x"5B",x"20",x"20",x"5D",x"20",x"20",x"42",x"2E",x"20", -- 3570-357F
  x"53",x"50",x"4D",x"45",x"52",x"4B",x"20",x"5B",x"20",x"5D",x"20",x"4F",x"42",x"4A",x"2B",x"30", -- 3580-358F
  x"20",x"4F",x"42",x"4A",x"44",x"55",x"4D",x"50",x"20",x"4F",x"42",x"4A",x"5F",x"53",x"54",x"52", -- 3590-359F
  x"55",x"43",x"54",x"5F",x"43",x"4F",x"50",x"59",x"20",x"53",x"49",x"5A",x"45",x"20",x"41",x"4D", -- 35A0-35AF
  x"45",x"52",x"4B",x"20",x"41",x"43",x"42",x"49",x"54",x"20",x"41",x"44",x"42",x"49",x"54",x"20", -- 35B0-35BF
  x"41",x"44",x"45",x"42",x"55",x"47",x"31",x"20",x"41",x"44",x"45",x"42",x"55",x"47",x"31",x"20", -- 35C0-35CF
  x"20",x"41",x"44",x"45",x"42",x"55",x"47",x"32",x"20",x"41",x"44",x"45",x"42",x"55",x"47",x"32", -- 35D0-35DF
  x"20",x"20",x"5B",x"41",x"2A",x"78",x"2D",x"59",x"2A",x"5A",x"5D",x"2F",x"67",x"78",x"20",x"49", -- 35E0-35EF
  x"4E",x"56",x"45",x"52",x"54",x"49",x"45",x"52",x"45",x"4E",x"20",x"56",x"41",x"4E",x"44",x"45", -- 35F0-35FF
  x"52",x"4D",x"4F",x"4E",x"44",x"45",x"4D",x"41",x"54",x"52",x"49",x"58",x"20",x"56",x"4C",x"49", -- 3600-360F
  x"53",x"54",x"20",x"57",x"4C",x"49",x"53",x"54",x"20",x"46",x"4F",x"52",x"47",x"45",x"54",x"20", -- 3610-361F
  x"6E",x"69",x"63",x"68",x"74",x"20",x"67",x"65",x"66",x"75",x"6E",x"64",x"65",x"6E",x"20",x"20", -- 3620-362F
  x"46",x"45",x"48",x"4C",x"45",x"52",x"54",x"45",x"58",x"54",x"20",x"44",x"69",x"76",x"69",x"73", -- 3630-363F
  x"69",x"6F",x"6E",x"20",x"64",x"75",x"72",x"63",x"68",x"20",x"4E",x"75",x"6C",x"6C",x"20",x"57", -- 3640-364F
  x"6F",x"72",x"74",x"20",x"6E",x"69",x"63",x"68",x"74",x"20",x"64",x"65",x"66",x"69",x"6E",x"69", -- 3650-365F
  x"65",x"72",x"74",x"20",x"45",x"69",x"6E",x"67",x"61",x"62",x"65",x"7A",x"65",x"69",x"6C",x"65", -- 3660-366F
  x"20",x"7A",x"75",x"20",x"6C",x"61",x"6E",x"67",x"20",x"53",x"74",x"72",x"75",x"6B",x"74",x"75", -- 3670-367F
  x"72",x"66",x"65",x"68",x"6C",x"65",x"72",x"20",x"69",x"6E",x"20",x"49",x"46",x"20",x"45",x"4E", -- 3680-368F
  x"44",x"5F",x"49",x"46",x"20",x"42",x"45",x"47",x"49",x"4E",x"20",x"55",x"4E",x"54",x"49",x"4C", -- 3690-369F
  x"20",x"44",x"4F",x"20",x"4C",x"4F",x"4F",x"50",x"20",x"20",x"6E",x"65",x"67",x"61",x"74",x"69", -- 36A0-36AF
  x"76",x"65",x"72",x"20",x"45",x"78",x"70",x"6F",x"6E",x"65",x"6E",x"74",x"20",x"5A",x"61",x"68", -- 36B0-36BF
  x"6C",x"65",x"6E",x"73",x"70",x"65",x"69",x"63",x"68",x"65",x"72",x"20",x"76",x"6F",x"6C",x"6C", -- 36C0-36CF
  x"20",x"67",x"72",x"6F",x"C3",x"9F",x"65",x"20",x"67",x"61",x"6E",x"7A",x"65",x"20",x"5A",x"61", -- 36D0-36DF
  x"68",x"6C",x"65",x"6E",x"20",x"6B",x"6F",x"6D",x"70",x"69",x"6C",x"69",x"65",x"72",x"65",x"6E", -- 36E0-36EF
  x"20",x"67",x"65",x"68",x"74",x"20",x"6D",x"6F",x"6D",x"65",x"6E",x"74",x"61",x"6E",x"20",x"6E", -- 36F0-36FF
  x"69",x"63",x"68",x"74",x"2E",x"20",x"53",x"54",x"52",x"47",x"3A",x"20",x"5E",x"47",x"20",x"2F", -- 3700-370F
  x"31",x"78",x"50",x"49",x"45",x"50",x"2F",x"20",x"5E",x"46",x"20",x"51",x"55",x"49",x"54",x"20", -- 3710-371F
  x"5E",x"41",x"20",x"41",x"6E",x"67",x"65",x"68",x"61",x"6C",x"74",x"65",x"6E",x"20",x"66",x"C3", -- 3720-372F
  x"BC",x"72",x"20",x"67",x"65",x"6E",x"61",x"75",x"20",x"65",x"69",x"6E",x"65",x"20",x"45",x"69", -- 3730-373F
  x"6E",x"67",x"61",x"62",x"65",x"7A",x"65",x"69",x"6C",x"65",x"3A",x"20",x"20",x"6F",x"6B",x"20", -- 3740-374F
  x"51",x"55",x"45",x"52",x"59",x"20",x"28",x"2A",x"52",x"45",x"4D",x"2A",x"29",x"20",x"2F",x"6F", -- 3750-375F
  x"6B",x"3E",x"20",x"28",x"2A",x"45",x"4E",x"44",x"2A",x"29",x"20",x"6F",x"6B",x"3E",x"20",x"48", -- 3760-376F
  x"45",x"58",x"20",x"44",x"45",x"43",x"49",x"4D",x"41",x"4C",x"20",x"3F",x"20",x"32",x"40",x"20", -- 3770-377F
  x"32",x"21",x"20",x"32",x"3F",x"20",x"52",x"41",x"4D",x"50",x"33",x"20",x"52",x"41",x"4D",x"42", -- 3780-378F
  x"55",x"46",x"20",x"54",x"4C",x"49",x"53",x"54",x"45",x"20",x"54",x"4C",x"49",x"53",x"54",x"45", -- 3790-379F
  x"4E",x"5A",x"45",x"49",x"47",x"45",x"52",x"20",x"54",x"4C",x"49",x"53",x"54",x"59",x"20",x"52", -- 37A0-37AF
  x"45",x"4D",x"4F",x"50",x"46",x"41",x"20",x"53",x"54",x"41",x"54",x"4D",x"45",x"52",x"4B",x"20", -- 37B0-37BF
  x"45",x"58",x"58",x"49",x"55",x"48",x"52",x"20",x"45",x"58",x"58",x"49",x"20",x"45",x"4E",x"54", -- 37C0-37CF
  x"46",x"45",x"52",x"4E",x"45",x"20",x"42",x"45",x"46",x"45",x"53",x"54",x"49",x"47",x"45",x"20", -- 37D0-37DF
  x"4C",x"49",x"4E",x"4B",x"53",x"2D",x"41",x"42",x"47",x"45",x"53",x"43",x"48",x"49",x"43",x"4B", -- 37E0-37EF
  x"54",x"20",x"52",x"45",x"43",x"48",x"54",x"53",x"2D",x"41",x"42",x"47",x"45",x"53",x"43",x"48", -- 37F0-37FF
  x"49",x"43",x"4B",x"54",x"20",x"4C",x"49",x"4E",x"4B",x"53",x"2D",x"41",x"4E",x"47",x"45",x"4B", -- 3800-380F
  x"4F",x"4D",x"4D",x"45",x"4E",x"20",x"52",x"45",x"43",x"48",x"54",x"53",x"2D",x"41",x"4E",x"47", -- 3810-381F
  x"45",x"4B",x"4F",x"4D",x"4D",x"45",x"4E",x"20",x"4F",x"42",x"45",x"4E",x"2D",x"41",x"42",x"47", -- 3820-382F
  x"45",x"53",x"43",x"48",x"49",x"43",x"4B",x"54",x"20",x"55",x"4E",x"54",x"45",x"4E",x"2D",x"41", -- 3830-383F
  x"42",x"47",x"45",x"53",x"43",x"48",x"49",x"43",x"4B",x"54",x"20",x"4F",x"42",x"45",x"4E",x"2D", -- 3840-384F
  x"41",x"4E",x"47",x"45",x"4B",x"4F",x"4D",x"4D",x"45",x"4E",x"20",x"55",x"4E",x"54",x"45",x"4E", -- 3850-385F
  x"2D",x"41",x"4E",x"47",x"45",x"4B",x"4F",x"4D",x"4D",x"45",x"4E",x"20",x"52",x"45",x"43",x"48", -- 3860-386F
  x"54",x"53",x"2D",x"42",x"59",x"54",x"45",x"53",x"20",x"55",x"4E",x"54",x"45",x"4E",x"2D",x"42", -- 3870-387F
  x"59",x"54",x"45",x"53",x"20",x"4C",x"49",x"4E",x"4B",x"53",x"2D",x"42",x"59",x"54",x"45",x"53", -- 3880-388F
  x"20",x"4F",x"42",x"45",x"4E",x"2D",x"42",x"59",x"54",x"45",x"53",x"20",x"49",x"41",x"4D",x"31", -- 3890-389F
  x"4A",x"20",x"49",x"41",x"4D",x"31",x"4B",x"20",x"49",x"41",x"4D",x"32",x"4A",x"20",x"49",x"41", -- 38A0-38AF
  x"4D",x"32",x"4B",x"20",x"4E",x"4A",x"20",x"4E",x"4B",x"20",x"4C",x"49",x"4E",x"4B",x"53",x"2D", -- 38B0-38BF
  x"4D",x"45",x"52",x"4B",x"20",x"4F",x"42",x"45",x"4E",x"2D",x"4D",x"45",x"52",x"4B",x"20",x"52", -- 38C0-38CF
  x"45",x"43",x"48",x"54",x"53",x"2D",x"4D",x"45",x"52",x"4B",x"20",x"55",x"4E",x"54",x"45",x"4E", -- 38D0-38DF
  x"2D",x"4D",x"45",x"52",x"4B",x"20",x"4A",x"4B",x"5F",x"41",x"55",x"53",x"47",x"45",x"42",x"20", -- 38E0-38EF
  x"52",x"2D",x"41",x"42",x"53",x"43",x"48",x"49",x"43",x"4B",x"45",x"4E",x"20",x"72",x"5F",x"77", -- 38F0-38FF
  x"61",x"72",x"74",x"20",x"20",x"55",x"2D",x"41",x"42",x"53",x"43",x"48",x"49",x"43",x"4B",x"45", -- 3900-390F
  x"4E",x"20",x"75",x"5F",x"77",x"61",x"72",x"74",x"20",x"20",x"41",x"42",x"53",x"43",x"48",x"49", -- 3910-391F
  x"43",x"4B",x"45",x"4E",x"20",x"41",x"42",x"57",x"41",x"52",x"54",x"20",x"4A",x"4B",x"2D",x"50", -- 3920-392F
  x"52",x"4F",x"43",x"20",x"3A",x"4B",x"20",x"20",x"4B",x"3A",x"20",x"20",x"42",x"5F",x"41",x"55", -- 3930-393F
  x"53",x"4C",x"45",x"53",x"20",x"42",x"5F",x"41",x"55",x"53",x"47",x"45",x"42",x"20",x"42",x"5F", -- 3940-394F
  x"49",x"4E",x"54",x"45",x"52",x"50",x"20",x"4C",x"2D",x"41",x"55",x"53",x"4C",x"45",x"53",x"20", -- 3950-395F
  x"4F",x"2D",x"41",x"55",x"53",x"4C",x"45",x"53",x"20",x"4E",x"20",x"4E",x"4E",x"20",x"4E",x"49", -- 3960-396F
  x"20",x"4A",x"4C",x"4F",x"43",x"20",x"4B",x"4C",x"4F",x"43",x"20",x"47",x"58",x"4D",x"45",x"52", -- 3970-397F
  x"4B",x"20",x"4D",x"2F",x"20",x"4A",x"4C",x"4F",x"43",x"21",x"20",x"4B",x"4C",x"4F",x"43",x"21", -- 3980-398F
  x"20",x"59",x"43",x"4F",x"4C",x"20",x"58",x"59",x"42",x"49",x"54",x"20",x"58",x"59",x"4D",x"45", -- 3990-399F
  x"52",x"4B",x"20",x"5A",x"42",x"49",x"54",x"20",x"5A",x"4D",x"45",x"52",x"4B",x"20",x"41",x"58", -- 39A0-39AF
  x"59",x"5A",x"20",x"58",x"59",x"53",x"50",x"45",x"49",x"43",x"48",x"20",x"5A",x"53",x"50",x"45", -- 39B0-39BF
  x"49",x"43",x"48",x"20",x"4D",x"2E",x"20",x"42",x"41",x"4E",x"46",x"20",x"40",x"20",x"34",x"30", -- 39C0-39CF
  x"20",x"54",x"59",x"50",x"45",x"20",x"20",x"3F",x"3F",x"3F",x"20",x"46",x"45",x"48",x"4C",x"45", -- 39D0-39DF
  x"52",x"54",x"45",x"58",x"54",x"20",x"45",x"52",x"52",x"4F",x"52",x"20",x"2D",x"20",x"46",x"65", -- 39E0-39EF
  x"68",x"6C",x"65",x"72",x"20",x"4E",x"75",x"6D",x"6D",x"65",x"72",x"20",x"20",x"5A",x"4C",x"4F", -- 39F0-39FF
  x"53",x"20",x"5A",x"4C",x"4F",x"53",x"20",x"20",x"58",x"59",x"4C",x"4F",x"53",x"20",x"58",x"59", -- 3A00-3A0F
  x"4C",x"4F",x"53",x"20",x"20",x"44",x"52",x"4F",x"50",x"20",x"5A",x"4C",x"4F",x"53",x"20",x"20", -- 3A10-3A1F
  x"47",x"49",x"4E",x"56",x"20",x"47",x"49",x"4E",x"56",x"20",x"20",x"4E",x"20",x"21",x"20",x"20", -- 3A20-3A2F
  x"47",x"49",x"4E",x"56",x"20",x"20",x"6B",x"6C",x"4D",x"61",x"74",x"41",x"75",x"66",x"74",x"20", -- 3A30-3A3F
  x"44",x"52",x"4F",x"50",x"20",x"5B",x"20",x"5B",x"20",x"20",x"44",x"52",x"4F",x"50",x"20",x"5D", -- 3A40-3A4F
  x"20",x"5B",x"20",x"20",x"44",x"52",x"4F",x"50",x"20",x"5D",x"20",x"5D",x"20",x"20",x"49",x"4E", -- 3A50-3A5F
  x"56",x"45",x"52",x"54",x"49",x"45",x"52",x"45",x"5F",x"53",x"43",x"48",x"4E",x"45",x"4C",x"4C", -- 3A60-3A6F
  x"20",x"61",x"30",x"30",x"2B",x"64",x"20",x"61",x"30",x"30",x"2B",x"64",x"20",x"20",x"30",x"41", -- 3A70-3A7F
  x"4D",x"45",x"52",x"4B",x"21",x"20",x"5A",x"55",x"52",x"55",x"45",x"43",x"4B",x"53",x"43",x"48", -- 3A80-3A8F
  x"49",x"43",x"4B",x"45",x"4E",x"20",x"42",x"28",x"6A",x"2C",x"6B",x"29",x"40",x"20",x"41",x"55", -- 3A90-3A9F
  x"53",x"47",x"41",x"4E",x"47",x"53",x"4D",x"41",x"54",x"52",x"49",x"58",x"5F",x"4E",x"55",x"4C", -- 3AA0-3AAF
  x"4C",x"53",x"45",x"54",x"5A",x"45",x"4E",x"20",x"48",x"41",x"55",x"50",x"54",x"4E",x"45",x"4E", -- 3AB0-3ABF
  x"4E",x"45",x"52",x"20",x"41",x"6A",x"6B",x"21",x"20",x"41",x"28",x"6A",x"2C",x"6B",x"29",x"21", -- 3AC0-3ACF
  x"20",x"56",x"41",x"4E",x"44",x"45",x"52",x"4D",x"4F",x"4E",x"44",x"45",x"4D",x"41",x"54",x"52", -- 3AD0-3ADF
  x"49",x"58",x"5F",x"47",x"4C",x"45",x"49",x"43",x"48",x"5F",x"41",x"55",x"46",x"54",x"45",x"49", -- 3AE0-3AEF
  x"4C",x"45",x"4E",x"20",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00", -- 3AF0-3AFF

  others=>x"00");

-- Rückkehrstapel
type stapRAMTYPE is array(0 to 1024-1) of STD_LOGIC_VECTOR (15 downto 0);
shared variable stapR: stapRAMTYPE:=(

  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C00-2C0F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C10-2C1F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C20-2C2F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C30-2C3F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C40-2C4F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C50-2C5F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C60-2C6F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C70-2C7F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C80-2C8F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2C90-2C9F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2CA0-2CAF
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2CB0-2CBF
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2CC0-2CCF
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2CD0-2CDF
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2CE0-2CEF
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2CF0-2CFF
  x"0000",x"0000",x"0000",x"0000",x"0055",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D00-2D0F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D10-2D1F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D20-2D2F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D30-2D3F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D40-2D4F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D50-2D5F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D60-2D6F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D70-2D7F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D80-2D8F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2D90-2D9F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2DA0-2DAF
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2DB0-2DBF
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2DC0-2DCF
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2DD0-2DDF
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2DE0-2DEF
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2DF0-2DFF
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E00-2E0F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E10-2E1F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E20-2E2F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E30-2E3F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E40-2E4F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E50-2E5F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E60-2E6F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E70-2E7F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E80-2E8F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2E90-2E9F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2EA0-2EAF
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2EB0-2EBF
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2EC0-2ECF
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2ED0-2EDF
  x"1667",x"16D6",x"0000",x"0000",x"0000",x"0000",x"0008",x"0000",x"0002",x"1E4E",x"0000",x"0001",x"2F22",x"1E4F",x"0009",x"1D9D", -- 2EE0-2EEF
  x"0008",x"0000",x"0001",x"2F22",x"0000",x"0001",x"2F23",x"1C02",x"0008",x"3B0A",x"0001",x"0001",x"3B45",x"00BB",x"0001",x"FFFF", -- 2EF0-2EFF
  x"0000",x"0000",x"3000",x"3E97",x"3E97",x"0000",x"3AF4",x"1B5D",x"0010",x"3B00",x"3B00",x"3B0C",x"3B12",x"3B45",x"0000",x"1B5D", -- 2F00-2F0F
  x"0000",x"1B22",x"3000",x"3AF4",x"0020",x"0020",x"0000",x"2D00",x"0000",x"1282",x"0000",x"0000",x"0000",x"0000",x"1277",x"126D", -- 2F10-2F1F
  x"2F47",x"0000",x"0000",x"1C00",x"1C00",x"2000",x"0001",x"0000",x"1C00",x"1C00",x"0000",x"FFD9",x"0000",x"0000",x"2EE0",x"2EE2", -- 2F20-2F2F
  x"16D6",x"0000",x"0000",x"FFFF",x"FFFF",x"FFFF",x"FFFF",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F30-2F3F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F40-2F4F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F50-2F5F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F60-2F6F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F70-2F7F
  x"2D00",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F80-2F8F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2F90-2F9F
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2FA0-2FAF
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2FB0-2FBF
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000", -- 2FC0-2FCF
  x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0301",x"0301",x"0301",x"0301",x"0301",x"0301",x"0301",x"0301", -- 2FD0-2FDF
  x"0301",x"0301",x"0301",x"0301",x"0446",x"02D5",x"02CD",x"02A3",x"02A3",x"02A3",x"02AB",x"02D6",x"02D6",x"0651",x"02D6",x"02D6", -- 2FE0-2FEF
  x"02D6",x"0624",x"02D6",x"02D6",x"031F",x"0345",x"01F6",x"029C",x"0812",x"FFFF",x"06EE",x"3B05",x"3B06",x"3B00",x"3B00",x"0738", -- 2FF0-2FFF

  others=>x"0000");

-- Datenspeicher 4000H-5FFFH
type DATRAMTYPE is array(0 to 8*1024-1) of STD_LOGIC_VECTOR (15 downto 0);
signal DatRAM: DATRAMTYPE:=(others=>x"0000");
-- RECHTS,UNTEN
type RUTYPE is array(0 to 1024-1) of STD_LOGIC_VECTOR (15 downto 0);
shared variable RechtsRAM: RUTYPE:=(others=>x"0000");
shared variable UntenRAM: RUTYPE:=(others=>x"0000");

--diese Funktion übernimmt von SP nur die beiden niedrigsten Bits
  function P(SP : integer) return integer is begin
--    return CONV_INTEGER(CONV_UNSIGNED(SP,2));
    return SP mod 4;
    end;

-- alles Signale um die Stapel-RAM's zu machen.
signal HOLE_VOM_STAPEL,STORE_ZUM_STAPEL,ADRESSE_ZUM_STAPEL: REG;
signal WE_ZUM_STAPEL: STD_LOGIC_VECTOR (3 downto 0);
type STAPELTYPE is array(0 to 31) of STD_LOGIC_VECTOR (15 downto 0);
signal stap1,stap2,stap3,stap0: STAPELTYPE:=(others=>x"0000");
-- Rueckkehrstapel
signal RPC,RPCC: STD_LOGIC_VECTOR (15 downto 0);
signal RP: STD_LOGIC_VECTOR (15 downto 0):=x"3000";
signal RW: STD_LOGIC;
-- kompletten Speicher anschliessen
signal PC_ZUM_ProgRAM,PD_VOM_ProgRAM: STD_LOGIC_VECTOR (15 downto 0);
signal STORE_ZUM_RAM,EXFET,ADRESSE_ZUM_RAM: STD_LOGIC_VECTOR (15 downto 0);
signal FETCH_VOM_ProgRAM,FETCH_VOM_ByteRAM,FETCH_VOM_DatRAM,FETCH_VOM_stapR: STD_LOGIC_VECTOR (15 downto 0);
signal WE_ZUM_RAM,WE_ZUM_ProgRAM,WE_ZUM_ByteRAM,WE_ZUM_DatRAM,WE_ZUM_stapR: STD_LOGIC;
-- fuer EMIT-Ausgabe
signal EMIT_ABGESCHICKT_LOCAL,EMIT_ANGEKOMMEN_RUHEND,XOFF_INPUT_L: STD_LOGIC:='0';
signal KEY_ANGEKOMMEN_LOCAL,KEY_ABGESCHICKT_RUHEND,KEY_ABGESCHICKT_MERK: STD_LOGIC:='0';
signal KEY_BYTE_RUHEND: STD_LOGIC_VECTOR (7 downto 0);
-- fuer LINKS-RECHTS-OBEN-UNTEN
signal LINKS_ABGESCHICKT_RUHEND,RECHTS_ANGEKOMMEN_RUHEND: STD_LOGIC:='0';
signal WE_ZUM_RechtsRAM: STD_LOGIC:='0';
signal OBEN_ABGESCHICKT_RUHEND,UNTEN_ANGEKOMMEN_RUHEND: STD_LOGIC:='0';
signal WE_ZUM_UntenRAM: STD_LOGIC:='0';


begin

process begin wait until (CLK_I'event and CLK_I='1'); --ruhende Eingangsdaten für FortyForthprocessor
  EMIT_ANGEKOMMEN_RUHEND<=EMIT_ANGEKOMMEN;
  KEY_BYTE_RUHEND<=KEY_BYTE;
  KEY_ABGESCHICKT_RUHEND<=KEY_ABGESCHICKT;
  LINKS_ABGESCHICKT_RUHEND<=LINKS_ABGESCHICKT;
  RECHTS_ANGEKOMMEN_RUHEND<=RECHTS_ANGEKOMMEN;
  OBEN_ABGESCHICKT_RUHEND<=OBEN_ABGESCHICKT;
  UNTEN_ANGEKOMMEN_RUHEND<=UNTEN_ANGEKOMMEN;
  end process;
  

process -- FortyForthProcessor
variable PC,PD,ADR,DAT,DIST: STD_LOGIC_VECTOR (15 downto 0):=x"0000";
variable WE: STD_LOGIC;
variable SP: integer:=0;
variable R: REG:=(others=>x"0000");
-- Stapeleintraege benennen
variable A,B,C,D: STD_LOGIC_VECTOR (15 downto 0):=x"0000";
variable T: integer range 0 to 4;
variable W: STD_LOGIC_VECTOR (3 downto 0);
-- fuer Umstapeln 
variable STAK: STD_LOGIC_VECTOR (7 downto 0);
-- fuer Rechenoperationen mit Uebertrag
variable U: STD_LOGIC_VECTOR (31 downto 0);
-- fuer Division
variable UBIT: STD_LOGIC;
-- fuer Supermult
variable SUMME: STD_LOGIC_VECTOR (31 downto 0);

begin wait until (CLK_I'event and CLK_I='0'); PC_SIM<=PC;--Simulation
  -- ob ein KEY aingetroffen ist --
  if KEY_ABGESCHICKT_MERK/=KEY_ABGESCHICKT_RUHEND then 
    KEY_ABGESCHICKT_MERK<=KEY_ABGESCHICKT_RUHEND;
    PD:=x"4012";
    PC:=PC;
    else
      PD:=PD_VOM_ProgRAM;
      PC:=PC+1;
      end if;                                           -- Simulation --
  WE:='0';                                              PD_SIM<=PD;
  DIST:=PD(11)&PD(11)&PD(11)&PD(11)&PD(11 downto 0);    SP_SIM<=CONV_STD_LOGIC_VECTOR(SP,16);
  -- oberste 4 Stapeleintraege entnehmen
  R:=HOLE_VOM_STAPEL;                                   -- Simulation --
  A:=R(P(SP-1));                                        A_SIM<=A;
  B:=R(P(SP-2));                                        B_SIM<=B;
  C:=R(P(SP-3));                                        C_SIM<=C;
  D:=R(P(SP-4));                                        D_SIM<=D;
  T:=0;
  -- Rueckkehrstapel
  RW<='0';
 
  if PD(15 downto 13)="010" then                 -- 4000-5FFF Unterprogrammaufruf
    RPC<=PC;PC:=PD and x"3FFF";RP<=RP-1;RW<='1';
    elsif PD(15 downto 12)=x"8" then PC:=PC+DIST;-- 8000-8FFF relativer Sprung
    elsif PD(15 downto 12)=x"9" then             -- 9000-9FFF bedingter relativer Sprung
      if A=x"0000" then PC:=PC+DIST; end if; SP:=SP-1;
    elsif PD=x"A003" then PC:=RPCC;RP<=RP+1;     -- ; Rückkehr aus Unterprogramm
    elsif PD=x"A00D" then -- 0= Vergleich ob gleich Null
      if A=x"0000" then A:=x"FFFF"; 
        else A:=x"0000"; end if;
      T:=1;
    elsif PD=x"A00F" then -- 0< Vergleich ob kleiner Null
      if A>=x"8000" then A:=x"FFFF";
        else A:=x"0000"; end if;
      T:=1;
    elsif PD=x"A000" then -- MINUS Vorzeichen wechseln
      A:=(not A)+1;
      T:=1;
    elsif PD=x"A00B" then -- NOT Bitweises Komplement
      A:=not A;
      T:=1;
    elsif PD=x"A008" then -- AND Bitweises Und
      A:=B and A; 
      T:=1;
      SP:=SP-1;
    elsif PD=x"A00E" then -- OR Bitweises Oder
      A:=B or A; 
      T:=1;
      SP:=SP-1;
    elsif PD=x"A007" then -- + Addition
      A:=B+A; 
      T:=1;
      SP:=SP-1;
    elsif PD=x"A001" then -- U+ Addition mit Übertrag
      U:=(x"0000"&C)+(x"0000"&B)+(x"0000"&A);
      B:=U(31 downto 16);
      A:=U(15 downto 0);
      T:=2;
      SP:=SP-1;
    elsif PD=x"A002" then -- U* Multiplikation mit Übertrag
      U:=(x"0000"&C)+B*A;
      B:=U(31 downto 16);
      A:=U(15 downto 0);
      T:=2;
      SP:=SP-1;
    elsif PD=x"A005" then -- EMIT Zeichen ausgeben
      if (EMIT_ABGESCHICKT_LOCAL=EMIT_ANGEKOMMEN_RUHEND) and XOFF_INPUT_L='0' then
        EMIT_BYTE<=A(7 downto 0);
        EMIT_ABGESCHICKT_LOCAL<=not EMIT_ANGEKOMMEN_RUHEND;
        T:=0;
        SP:=SP-1;
        else PC:=PC-1; end if; -- warten
    elsif PD=x"A009" then -- STORE Speicheradresse beschreiben
      case A is
        when x"2800" => KEY_ANGEKOMMEN_LOCAL<=not KEY_ANGEKOMMEN_LOCAL;
        when x"2801" => SP:=CONV_INTEGER(B);
        when x"2802" => RP<=B;
        when x"2803" => PC:=B;
        when x"2804" => RECHTS_ABGESCHICKT<=B(0);
        when x"2805" => LINKS_ANGEKOMMEN<=B(0);
        when x"2806" => UNTEN_ABGESCHICKT<=B(0);
        when x"2807" => OBEN_ANGEKOMMEN<=B(0);
        when others => ADR:=A;DAT:=B;WE:='1' ;
        end case;
      T:=0;
      SP:=SP-2;
    elsif PD=x"A00A" then -- FETCH Speicheradresse lesen
      case A is
        when x"2800" => A:=x"00"&KEY_BYTE_RUHEND;
        when x"2801" => A:=CONV_STD_LOGIC_VECTOR(SP-1,16);
        when x"2802" => A:=RP;
        when x"2803" => A:=PC;
        when x"2804" => A:="000000000000000"&LINKS_ABGESCHICKT_RUHEND;
        when x"2805" => A:="000000000000000"&RECHTS_ANGEKOMMEN_RUHEND;
        when x"2806" => A:="000000000000000"&OBEN_ABGESCHICKT_RUHEND;
        when x"2807" => A:="000000000000000"&UNTEN_ANGEKOMMEN_RUHEND;
        when others => A:=EXFET;
        end case;
      T:=1;
    elsif PD=x"A014" then -- DI32 DIVISION_MIT_REST 32B/16B=16R/16Q
      UBIT:=C(15);
      C:=C(14 downto 0)&B(15);
      B:=B(14 downto 0)&'0';
      if (UBIT&C)>=('0'&A) then
        C:=C-A;
        B(0):='1';
        end if;
      T:=3;
    elsif PD=x"A017" then -- MULT_I
      --     D    C    B    A        stapR
      --     c    ü   adr1 adr2      i
      -- c   ü   erg1 adr2 adr1      i-1
      SUMME:=(D*EXFET)+(x"0000"&C);
      C:=A;A:=B;B:=C;
      D:=SUMME(31 downto 16); 
      C:=SUMME(15 downto 0);
      RPC<=RPCC-1; RW<='1';
      T:=4; SP:=SP+1;
    elsif PD=x"A018" then -- MULT_II
      --     D    C     B      A         stapR
      -- c   ü1  erg1   adr2   adr1      i-1
      -- c   ü2  adr1+1 adr2+1 i-1       i-1
      SUMME:=(D&C)+(x"0000"&EXFET);
      D:=SUMME(31 downto 16); 
      DAT:=SUMME(15 downto 0);
      ADR:=A;
      WE:='1';
      C:=A+1;
      B:=B+1;
      if RPCC=x"0000" then A:=x"FFFF"; else A:=x"0000"; end if;
      T:=4;
    elsif PD(15 downto 12)=x"B" then           -- B000-BFFF Umstapeln
      STAK:="00000000";
      if PD(7)='1' then STAK:=STAK(5 downto 0)&"11"; T:=T+1; end if;
      if PD(6)='1' then STAK:=STAK(5 downto 0)&"10"; T:=T+1; end if;
      if PD(5)='1' then STAK:=STAK(5 downto 0)&"01"; T:=T+1; end if;
      if PD(4)='1' then STAK:=STAK(5 downto 0)&"00"; T:=T+1; end if;
      if PD(3)='1' then STAK:=STAK(5 downto 0)&"11"; T:=T+1; end if;
      if PD(2)='1' then STAK:=STAK(5 downto 0)&"10"; T:=T+1; end if;
      if PD(1)='1' then STAK:=STAK(5 downto 0)&"01"; T:=T+1; end if;
      if PD(0)='1' then STAK:=STAK(5 downto 0)&"00"; T:=T+1; end if;
      A:=R(P(SP-1-CONV_INTEGER(STAK(1 downto 0))));
      B:=R(P(SP-1-CONV_INTEGER(STAK(3 downto 2))));
      C:=R(P(SP-1-CONV_INTEGER(STAK(5 downto 4))));
      D:=R(P(SP-1-CONV_INTEGER(STAK(7 downto 6))));
      SP:=SP+CONV_INTEGER(PD(11 downto 8))-4;
    else A:=PD; SP:=SP+1; T:=1; end if;                    -- LIT
    
  -- oberste T Stapeleintraege zurückspeichern
  W:="0000";
  if T/=0 then R(P(SP-1)):=A; W(P(SP-1)):='1';
    if T/=1 then R(P(SP-2)):=B; W(P(SP-2)):='1';
      if T/=2 then R(P(SP-3)):=C; W(P(SP-3)):='1';
        if T/=3 then R(P(SP-4)):=D; W(P(SP-4)):='1';
          end if; end if; end if; end if;
  -- Ausgabeadresse zum StapRAM zusammenbasteln
  ADRESSE_ZUM_STAPEL(0)<=CONV_STD_LOGIC_VECTOR(SP-1,16);
  ADRESSE_ZUM_STAPEL(1)<=CONV_STD_LOGIC_VECTOR(SP-2,16);
  ADRESSE_ZUM_STAPEL(2)<=CONV_STD_LOGIC_VECTOR(SP-3,16);
  ADRESSE_ZUM_STAPEL(3)<=CONV_STD_LOGIC_VECTOR(SP-4,16);
  STORE_ZUM_STAPEL<=R;
  WE_ZUM_STAPEL<=W;
  -- ADR, DAT, WE, PC
  if WE='1' then ADRESSE_ZUM_RAM<=ADR; else ADRESSE_ZUM_RAM<=R(P(SP-1)); end if;
  STORE_ZUM_RAM<=DAT;
  WE_ZUM_RAM<=WE;
  PC_ZUM_ProgRAM<=PC;
  end process;

ADR_O<=ADRESSE_ZUM_RAM;
DAT_O<=STORE_ZUM_RAM;
WE_O<=WE_ZUM_RAM;
EMIT_ABGESCHICKT<=EMIT_ABGESCHICKT_LOCAL;
KEY_ANGEKOMMEN<=KEY_ANGEKOMMEN_LOCAL;
LINKS_ADR<=ADRESSE_ZUM_RAM;
OBEN_ADR<=ADRESSE_ZUM_RAM;

-- hier werden die Lesedaten der unterschiedlichen Speicher zusammengefuehrt
EXFET<=FETCH_VOM_ProgRAM when ADRESSE_ZUM_RAM(15 downto 13)="000" else
       FETCH_VOM_stapR when ADRESSE_ZUM_RAM(15 downto 10)="001011" else
       LINKS_DAT when ADRESSE_ZUM_RAM(15 downto 10)="011110" else
       OBEN_DAT when ADRESSE_ZUM_RAM(15 downto 10)="011111" else
       x"00"&FETCH_VOM_ByteRAM(7 downto 0) when ADRESSE_ZUM_RAM(15 downto 12)="0011" else
       FETCH_VOM_DatRAM when ADRESSE_ZUM_RAM(15 downto 13)="010" else
       DAT_I;

-- hier wird WE auf die unterschiedlichen Speicher aufgeteilt
WE_ZUM_ProgRAM<=WE_ZUM_RAM when ADRESSE_ZUM_RAM(15 downto 13)="000" else '0';
WE_ZUM_RechtsRAM<=WE_ZUM_RAM when ADRESSE_ZUM_RAM(15 downto 10)="011110" else '0';
WE_ZUM_UntenRAM<=WE_ZUM_RAM when ADRESSE_ZUM_RAM(15 downto 10)="011111" else '0';
WE_ZUM_stapR  <=WE_ZUM_RAM when ADRESSE_ZUM_RAM(15 downto 10)="001011" else '0';
WE_ZUM_ByteRAM<=WE_ZUM_RAM when ADRESSE_ZUM_RAM(15 downto 12)="0011" else '0';
WE_ZUM_DatRAM<=WE_ZUM_RAM when ADRESSE_ZUM_RAM(15 downto 13)="010" else '0';


process -- Programmspeicher 0000H-1FFFH,
begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_ProgRAM='1' then 
    ProgRAM(CONV_INTEGER(ADRESSE_ZUM_RAM(12 downto 0)))<=STORE_ZUM_RAM; 
    FETCH_VOM_ProgRAM<=STORE_ZUM_RAM; 
	  else
      FETCH_VOM_ProgRAM<=ProgRAM(CONV_INTEGER(ADRESSE_ZUM_RAM(12 downto 0)));
      end if;
  PD_VOM_ProgRAM<=ProgRAM(CONV_INTEGER(PC_ZUM_ProgRAM(12 downto 0)));
  end process;

process -- Textspeicher 3000H-3FFFH
begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_ByteRAM='1' then 
    ByteRAM(CONV_INTEGER(ADRESSE_ZUM_RAM(11 downto 0)))<=STORE_ZUM_RAM(7 downto 0); 
    FETCH_VOM_ByteRAM<=STORE_ZUM_RAM; 
	 else
      FETCH_VOM_ByteRAM<=x"00"&ByteRAM(CONV_INTEGER(ADRESSE_ZUM_RAM(11 downto 0)));
      end if;
  end process;

process --Rueckkehrstapel, TRUE_DUAL_PORT
begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_StapR='1' then 
    stapR(CONV_INTEGER(ADRESSE_ZUM_RAM(9 downto 0))):=STORE_ZUM_RAM; 
    end if;
  FETCH_VOM_stapR<=stapR(CONV_INTEGER(ADRESSE_ZUM_RAM(9 downto 0)));
  end process;
process begin wait until (CLK_I'event and CLK_I='1');
  if RW='1' then
    stapR(CONV_INTEGER(RP(9 downto 0))):=RPC;
    RPCC<=RPC;
     else
      RPCC<=stapR(CONV_INTEGER(RP(9 downto 0)));
    end if;
  end process;

process -- Datenpeicher 4000H-5FFFH,
begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_DatRAM='1' then 
    DatRAM(CONV_INTEGER(ADRESSE_ZUM_RAM(12 downto 0)))<=STORE_ZUM_RAM; 
    FETCH_VOM_DatRAM<=STORE_ZUM_RAM; 
	  else
      FETCH_VOM_DatRAM<=DatRAM(CONV_INTEGER(ADRESSE_ZUM_RAM(12 downto 0)));
      end if;
  end process;

--StapelRAM:
process begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_STAPEL(0)='1' then
    stap0(CONV_INTEGER(ADRESSE_ZUM_STAPEL(0)(6 downto 2)))<=STORE_ZUM_STAPEL(0);
    HOLE_VOM_STAPEL(0)<=STORE_ZUM_STAPEL(0);
     else
      HOLE_VOM_STAPEL(0)<=stap0(CONV_INTEGER(ADRESSE_ZUM_STAPEL(0)(6 downto 2)));
    end if;
  end process;
process begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_STAPEL(1)='1' then
    stap1(CONV_INTEGER(ADRESSE_ZUM_STAPEL(1)(6 downto 2)))<=STORE_ZUM_STAPEL(1);
    HOLE_VOM_STAPEL(1)<=STORE_ZUM_STAPEL(1);
     else
      HOLE_VOM_STAPEL(1)<=stap1(CONV_INTEGER(ADRESSE_ZUM_STAPEL(1)(6 downto 2)));
    end if;
  end process;
process begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_STAPEL(2)='1' then
    stap2(CONV_INTEGER(ADRESSE_ZUM_STAPEL(2)(6 downto 2)))<=STORE_ZUM_STAPEL(2);
    HOLE_VOM_STAPEL(2)<=STORE_ZUM_STAPEL(2);
     else
      HOLE_VOM_STAPEL(2)<=stap2(CONV_INTEGER(ADRESSE_ZUM_STAPEL(2)(6 downto 2)));
    end if;
  end process;
process begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_STAPEL(3)='1' then
    stap3(CONV_INTEGER(ADRESSE_ZUM_STAPEL(3)(6 downto 2)))<=STORE_ZUM_STAPEL(3);
    HOLE_VOM_STAPEL(3)<=STORE_ZUM_STAPEL(3);
     else
      HOLE_VOM_STAPEL(3)<=stap3(CONV_INTEGER(ADRESSE_ZUM_STAPEL(3)(6 downto 2)));
    end if;
  end process;

process --RechtsRAM --DUAL-PORT
begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_RechtsRAM='1' then 
    RechtsRAM(CONV_INTEGER(ADRESSE_ZUM_RAM(9 downto 0))):=STORE_ZUM_RAM; 
    end if;
  --FETCH_VOM_stapR<=stapR(CONV_INTEGER(ADRESSE_ZUM_RAM(9 downto 0)));
  end process;
process begin wait until (CLK_I'event and CLK_I='1');
  if false then
    --stapR(CONV_INTEGER(RP(9 downto 0))):=RPC;
    --RPCC<=RPC;
     else
      RECHTS_DAT<=RechtsRAM(CONV_INTEGER(RECHTS_ADR(9 downto 0)));
    end if;
  end process;

process --UntenRAM --DUAL-PORT
begin wait until (CLK_I'event and CLK_I='1');
  if WE_ZUM_UntenRAM='1' then 
    UntenRAM(CONV_INTEGER(ADRESSE_ZUM_RAM(9 downto 0))):=STORE_ZUM_RAM; 
    end if;
  --FETCH_VOM_stapR<=stapR(CONV_INTEGER(ADRESSE_ZUM_RAM(9 downto 0)));
  end process;
process begin wait until (CLK_I'event and CLK_I='1');
  if false then
    --stapR(CONV_INTEGER(RP(9 downto 0))):=RPC;
    --RPCC<=RPC;
     else
      UNTEN_DAT<=UntenRAM(CONV_INTEGER(UNTEN_ADR(9 downto 0)));
    end if;
  end process;




end Step_12;
